LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY MBE IS
   PORT( 
      A : in std_logic_vector(31 DOWNTO 0);
      B : in std_logic_vector(31 DOWNTO 0); 
		M : out std_logic_vector(63 downto 0));

END MBE;

architecture behavior of MBE is

	component HA is 
		port (A: in std_logic; 	
				B: in std_logic;    
				S : out	std_logic; 	
				Cout : out	std_logic);    
	end component HA;
	
	component FA is 
		port (A: in std_logic; 	
				B: in std_logic; 	
				Cin: in std_logic;    
				S : out	std_logic; 	
				Cout : out	std_logic);    
	end component FA;
	
	component PP_gen is 
		port( A : in std_logic_vector(31 DOWNTO 0);   
				B : in std_logic_vector(31 DOWNTO 0);   
				PP0 : out std_logic_vector(32 downto 0);   
				PP1 : out std_logic_vector(32 downto 0);   
				PP2 : out std_logic_vector(32 downto 0);  
				PP3 : out std_logic_vector(32 downto 0);   
				PP4 : out std_logic_vector(32 downto 0);   
				PP5 : out std_logic_vector(32 downto 0);   
				PP6 : out std_logic_vector(32 downto 0);   
				PP7 : out std_logic_vector(32 downto 0);   
				PP8 : out std_logic_vector(32 downto 0);   
				PP9 : out std_logic_vector(32 downto 0);   
				PP10 : out std_logic_vector(32 downto 0);  
				PP11 : out std_logic_vector(32 downto 0);   
				PP12 : out std_logic_vector(32 downto 0);   
				PP13 : out std_logic_vector(32 downto 0);   
				PP14 : out std_logic_vector(32 downto 0);   
				PP15 : out std_logic_vector(32 downto 0);   
				PP16 : out std_logic_vector(31 downto 0));   
	end component PP_gen;
	
signal PP0 : std_logic_vector(32 downto 0);
signal PP1 : std_logic_vector(32 downto 0);
signal PP2 : std_logic_vector(32 downto 0);
signal PP3 : std_logic_vector(32 downto 0);
signal PP4 : std_logic_vector(32 downto 0);
signal PP5 : std_logic_vector(32 downto 0);
signal PP6 : std_logic_vector(32 downto 0);
signal PP7 : std_logic_vector(32 downto 0);
signal PP8 : std_logic_vector(32 downto 0);
signal PP9 : std_logic_vector(32 downto 0);
signal PP10 : std_logic_vector(32 downto 0);
signal PP11 : std_logic_vector(32 downto 0);
signal PP12 : std_logic_vector(32 downto 0);
signal PP13 : std_logic_vector(32 downto 0);
signal PP14 : std_logic_vector(32 downto 0);
signal PP15 : std_logic_vector(32 downto 0);
signal PP16 : std_logic_vector(31 downto 0);

signal PP0_neg : std_logic;
signal PP1_neg : std_logic;
signal PP2_neg : std_logic;
signal PP3_neg : std_logic;
signal PP4_neg : std_logic;
signal PP5_neg : std_logic;
signal PP6_neg : std_logic;
signal PP7_neg : std_logic;
signal PP8_neg : std_logic;
signal PP9_neg : std_logic;
signal PP10_neg: std_logic;
signal PP11_neg : std_logic;
signal PP12_neg : std_logic;
signal PP13_neg : std_logic;
signal PP14_neg : std_logic;
signal PP15_neg : std_logic;
--signal PP16_neg : std_logic;
	
signal HA1_l6_c24_S : std_logic;
signal HA1_l6_c24_Cout : std_logic;
signal HA1_l6_c25_S : std_logic;
signal HA1_l6_c25_Cout : std_logic;
signal FA1_l6_c26_S : std_logic;
signal FA1_l6_c26_Cout : std_logic;
signal HA1_l6_c26_S : std_logic;
signal HA1_l6_c26_Cout : std_logic;
signal FA1_l6_c27_S : std_logic;
signal FA1_l6_c27_Cout : std_logic;
signal HA1_l6_c27_S : std_logic;
signal HA1_l6_c27_Cout : std_logic;
signal FA1_l6_c28_S : std_logic;
signal FA1_l6_c28_Cout : std_logic;
signal FA2_l6_c28_S : std_logic;
signal FA2_l6_c28_Cout : std_logic;
signal HA1_l6_c28_S : std_logic;
signal HA1_l6_c28_Cout : std_logic;
signal FA1_l6_c29_S : std_logic;
signal FA1_l6_c29_Cout : std_logic;
signal FA2_l6_c29_S : std_logic;
signal FA2_l6_c29_Cout : std_logic;
signal HA1_l6_c29_S : std_logic;
signal HA1_l6_c29_Cout : std_logic;
signal FA1_l6_c30_S : std_logic;
signal FA1_l6_c30_Cout : std_logic;
signal FA2_l6_c30_S : std_logic;
signal FA2_l6_c30_Cout : std_logic;
signal FA3_l6_c30_S : std_logic;
signal FA3_l6_c30_Cout : std_logic;
signal HA1_l6_c30_S : std_logic;
signal HA1_l6_c30_Cout : std_logic;
signal FA1_l6_c31_S : std_logic;
signal FA1_l6_c31_Cout : std_logic;
signal FA2_l6_c31_S : std_logic;
signal FA2_l6_c31_Cout : std_logic;
signal FA3_l6_c31_S : std_logic;
signal FA3_l6_c31_Cout : std_logic;
signal HA1_l6_c31_S : std_logic;
signal HA1_l6_c31_Cout : std_logic;
signal FA1_l6_c32_S : std_logic;
signal FA1_l6_c32_Cout : std_logic;
signal FA2_l6_c32_S : std_logic;
signal FA2_l6_c32_Cout : std_logic;
signal FA3_l6_c32_S : std_logic;
signal FA3_l6_c32_Cout : std_logic;
signal FA4_l6_c32_S : std_logic;
signal FA4_l6_c32_Cout : std_logic;
signal FA1_l6_c33_S : std_logic;
signal FA1_l6_c33_Cout : std_logic;
signal FA2_l6_c33_S : std_logic;
signal FA2_l6_c33_Cout : std_logic;
signal FA3_l6_c33_S : std_logic;
signal FA3_l6_c33_Cout : std_logic;
signal FA4_l6_c33_S : std_logic;
signal FA4_l6_c33_Cout : std_logic;
signal FA1_l6_c34_S : std_logic;
signal FA1_l6_c34_Cout : std_logic;
signal FA2_l6_c34_S : std_logic;
signal FA2_l6_c34_Cout : std_logic;
signal FA3_l6_c34_S : std_logic;
signal FA3_l6_c34_Cout : std_logic;
signal FA4_l6_c34_S : std_logic;
signal FA4_l6_c34_Cout : std_logic;
signal FA1_l6_c35_S : std_logic;
signal FA1_l6_c35_Cout : std_logic;
signal FA2_l6_c35_S : std_logic;
signal FA2_l6_c35_Cout : std_logic;
signal FA3_l6_c35_S : std_logic;
signal FA3_l6_c35_Cout : std_logic;
signal FA4_l6_c35_S : std_logic;
signal FA4_l6_c35_Cout : std_logic;
signal FA1_l6_c36_S : std_logic;
signal FA1_l6_c36_Cout : std_logic;
signal FA2_l6_c36_S : std_logic;
signal FA2_l6_c36_Cout : std_logic;
signal FA3_l6_c36_S : std_logic;
signal FA3_l6_c36_Cout : std_logic;
signal HA1_l6_c36_S : std_logic;
signal HA1_l6_c36_Cout : std_logic;
signal FA1_l6_c37_S : std_logic;
signal FA1_l6_c37_Cout : std_logic;
signal FA2_l6_c37_S : std_logic;
signal FA2_l6_c37_Cout : std_logic;
signal FA3_l6_c37_S : std_logic;
signal FA3_l6_c37_Cout : std_logic;
signal FA1_l6_c38_S : std_logic;
signal FA1_l6_c38_Cout : std_logic;
signal FA2_l6_c38_S : std_logic;
signal FA2_l6_c38_Cout : std_logic;
signal HA1_l6_c38_S : std_logic;
signal HA1_l6_c38_Cout : std_logic;
signal FA1_l6_c39_S : std_logic;
signal FA1_l6_c39_Cout : std_logic;
signal FA2_l6_c39_S : std_logic;
signal FA2_l6_c39_Cout : std_logic;
signal FA1_l6_c40_S : std_logic;
signal FA1_l6_c40_Cout : std_logic;
signal HA1_l6_c40_S : std_logic;
signal HA1_l6_c40_Cout : std_logic;
signal FA1_l6_c41_S : std_logic;
signal FA1_l6_c41_Cout : std_logic;
signal HA1_l6_c42_S : std_logic;
signal HA1_l6_c42_Cout : std_logic;
signal HA1_l5_c16_S : std_logic;
signal HA1_l5_c16_Cout : std_logic;
signal HA1_l5_c17_S : std_logic;
signal HA1_l5_c17_Cout : std_logic;
signal FA1_l5_c18_S : std_logic;
signal FA1_l5_c18_Cout : std_logic;
signal HA1_l5_c18_S : std_logic;
signal HA1_l5_c18_Cout : std_logic;
signal FA1_l5_c19_S : std_logic;
signal FA1_l5_c19_Cout : std_logic;
signal HA1_l5_c19_S : std_logic;
signal HA1_l5_c19_Cout : std_logic;
signal FA1_l5_c20_S : std_logic;
signal FA1_l5_c20_Cout : std_logic;
signal FA2_l5_c20_S : std_logic;
signal FA2_l5_c20_Cout : std_logic;
signal HA1_l5_c20_S : std_logic;
signal HA1_l5_c20_Cout : std_logic;
signal FA1_l5_c21_S : std_logic;
signal FA1_l5_c21_Cout : std_logic;
signal FA2_l5_c21_S : std_logic;
signal FA2_l5_c21_Cout : std_logic;
signal HA1_l5_c21_S : std_logic;
signal HA1_l5_c21_Cout : std_logic;
signal FA1_l5_c22_S : std_logic;
signal FA1_l5_c22_Cout : std_logic;
signal FA2_l5_c22_S : std_logic;
signal FA2_l5_c22_Cout : std_logic;
signal FA3_l5_c22_S : std_logic;
signal FA3_l5_c22_Cout : std_logic;
signal HA1_l5_c22_S : std_logic;
signal HA1_l5_c22_Cout : std_logic;
signal FA1_l5_c23_S : std_logic;
signal FA1_l5_c23_Cout : std_logic;
signal FA2_l5_c23_S : std_logic;
signal FA2_l5_c23_Cout : std_logic;
signal FA3_l5_c23_S : std_logic;
signal FA3_l5_c23_Cout : std_logic;
signal HA1_l5_c23_S : std_logic;
signal HA1_l5_c23_Cout : std_logic;
signal FA1_l5_c24_S : std_logic;
signal FA1_l5_c24_Cout : std_logic;
signal FA2_l5_c24_S : std_logic;
signal FA2_l5_c24_Cout : std_logic;
signal FA3_l5_c24_S : std_logic;
signal FA3_l5_c24_Cout : std_logic;
signal FA4_l5_c24_S : std_logic;
signal FA4_l5_c24_Cout : std_logic;
signal FA1_l5_c25_S : std_logic;
signal FA1_l5_c25_Cout : std_logic;
signal FA2_l5_c25_S : std_logic;
signal FA2_l5_c25_Cout : std_logic;
signal FA3_l5_c25_S : std_logic;
signal FA3_l5_c25_Cout : std_logic;
signal FA4_l5_c25_S : std_logic;
signal FA4_l5_c25_Cout : std_logic;
signal FA1_l5_c26_S : std_logic;
signal FA1_l5_c26_Cout : std_logic;
signal FA2_l5_c26_S : std_logic;
signal FA2_l5_c26_Cout : std_logic;
signal FA3_l5_c26_S : std_logic;
signal FA3_l5_c26_Cout : std_logic;
signal FA4_l5_c26_S : std_logic;
signal FA4_l5_c26_Cout : std_logic;
signal FA1_l5_c27_S : std_logic;
signal FA1_l5_c27_Cout : std_logic;
signal FA2_l5_c27_S : std_logic;
signal FA2_l5_c27_Cout : std_logic;
signal FA3_l5_c27_S : std_logic;
signal FA3_l5_c27_Cout : std_logic;
signal FA4_l5_c27_S : std_logic;
signal FA4_l5_c27_Cout : std_logic;
signal FA1_l5_c28_S : std_logic;
signal FA1_l5_c28_Cout : std_logic;
signal FA2_l5_c28_S : std_logic;
signal FA2_l5_c28_Cout : std_logic;
signal FA3_l5_c28_S : std_logic;
signal FA3_l5_c28_Cout : std_logic;
signal FA4_l5_c28_S : std_logic;
signal FA4_l5_c28_Cout : std_logic;
signal FA1_l5_c29_S : std_logic;
signal FA1_l5_c29_Cout : std_logic;
signal FA2_l5_c29_S : std_logic;
signal FA2_l5_c29_Cout : std_logic;
signal FA3_l5_c29_S : std_logic;
signal FA3_l5_c29_Cout : std_logic;
signal FA4_l5_c29_S : std_logic;
signal FA4_l5_c29_Cout : std_logic;
signal FA1_l5_c30_S : std_logic;
signal FA1_l5_c30_Cout : std_logic;
signal FA2_l5_c30_S : std_logic;
signal FA2_l5_c30_Cout : std_logic;
signal FA3_l5_c30_S : std_logic;
signal FA3_l5_c30_Cout : std_logic;
signal FA4_l5_c30_S : std_logic;
signal FA4_l5_c30_Cout : std_logic;
signal FA1_l5_c31_S : std_logic;
signal FA1_l5_c31_Cout : std_logic;
signal FA2_l5_c31_S : std_logic;
signal FA2_l5_c31_Cout : std_logic;
signal FA3_l5_c31_S : std_logic;
signal FA3_l5_c31_Cout : std_logic;
signal FA4_l5_c31_S : std_logic;
signal FA4_l5_c31_Cout : std_logic;
signal FA1_l5_c32_S : std_logic;
signal FA1_l5_c32_Cout : std_logic;
signal FA2_l5_c32_S : std_logic;
signal FA2_l5_c32_Cout : std_logic;
signal FA3_l5_c32_S : std_logic;
signal FA3_l5_c32_Cout : std_logic;
signal FA4_l5_c32_S : std_logic;
signal FA4_l5_c32_Cout : std_logic;
signal FA1_l5_c33_S : std_logic;
signal FA1_l5_c33_Cout : std_logic;
signal FA2_l5_c33_S : std_logic;
signal FA2_l5_c33_Cout : std_logic;
signal FA3_l5_c33_S : std_logic;
signal FA3_l5_c33_Cout : std_logic;
signal FA4_l5_c33_S : std_logic;
signal FA4_l5_c33_Cout : std_logic;
signal FA1_l5_c34_S : std_logic;
signal FA1_l5_c34_Cout : std_logic;
signal FA2_l5_c34_S : std_logic;
signal FA2_l5_c34_Cout : std_logic;
signal FA3_l5_c34_S : std_logic;
signal FA3_l5_c34_Cout : std_logic;
signal FA4_l5_c34_S : std_logic;
signal FA4_l5_c34_Cout : std_logic;
signal FA1_l5_c35_S : std_logic;
signal FA1_l5_c35_Cout : std_logic;
signal FA2_l5_c35_S : std_logic;
signal FA2_l5_c35_Cout : std_logic;
signal FA3_l5_c35_S : std_logic;
signal FA3_l5_c35_Cout : std_logic;
signal FA4_l5_c35_S : std_logic;
signal FA4_l5_c35_Cout : std_logic;
signal FA1_l5_c36_S : std_logic;
signal FA1_l5_c36_Cout : std_logic;
signal FA2_l5_c36_S : std_logic;
signal FA2_l5_c36_Cout : std_logic;
signal FA3_l5_c36_S : std_logic;
signal FA3_l5_c36_Cout : std_logic;
signal FA4_l5_c36_S : std_logic;
signal FA4_l5_c36_Cout : std_logic;
signal FA1_l5_c37_S : std_logic;
signal FA1_l5_c37_Cout : std_logic;
signal FA2_l5_c37_S : std_logic;
signal FA2_l5_c37_Cout : std_logic;
signal FA3_l5_c37_S : std_logic;
signal FA3_l5_c37_Cout : std_logic;
signal FA4_l5_c37_S : std_logic;
signal FA4_l5_c37_Cout : std_logic;
signal FA1_l5_c38_S : std_logic;
signal FA1_l5_c38_Cout : std_logic;
signal FA2_l5_c38_S : std_logic;
signal FA2_l5_c38_Cout : std_logic;
signal FA3_l5_c38_S : std_logic;
signal FA3_l5_c38_Cout : std_logic;
signal FA4_l5_c38_S : std_logic;
signal FA4_l5_c38_Cout : std_logic;
signal FA1_l5_c39_S : std_logic;
signal FA1_l5_c39_Cout : std_logic;
signal FA2_l5_c39_S : std_logic;
signal FA2_l5_c39_Cout : std_logic;
signal FA3_l5_c39_S : std_logic;
signal FA3_l5_c39_Cout : std_logic;
signal FA4_l5_c39_S : std_logic;
signal FA4_l5_c39_Cout : std_logic;
signal FA1_l5_c40_S : std_logic;
signal FA1_l5_c40_Cout : std_logic;
signal FA2_l5_c40_S : std_logic;
signal FA2_l5_c40_Cout : std_logic;
signal FA3_l5_c40_S : std_logic;
signal FA3_l5_c40_Cout : std_logic;
signal FA4_l5_c40_S : std_logic;
signal FA4_l5_c40_Cout : std_logic;
signal FA1_l5_c41_S : std_logic;
signal FA1_l5_c41_Cout : std_logic;
signal FA2_l5_c41_S : std_logic;
signal FA2_l5_c41_Cout : std_logic;
signal FA3_l5_c41_S : std_logic;
signal FA3_l5_c41_Cout : std_logic;
signal FA4_l5_c41_S : std_logic;
signal FA4_l5_c41_Cout : std_logic;
signal FA1_l5_c42_S : std_logic;
signal FA1_l5_c42_Cout : std_logic;
signal FA2_l5_c42_S : std_logic;
signal FA2_l5_c42_Cout : std_logic;
signal FA3_l5_c42_S : std_logic;
signal FA3_l5_c42_Cout : std_logic;
signal FA4_l5_c42_S : std_logic;
signal FA4_l5_c42_Cout : std_logic;
signal FA1_l5_c43_S : std_logic;
signal FA1_l5_c43_Cout : std_logic;
signal FA2_l5_c43_S : std_logic;
signal FA2_l5_c43_Cout : std_logic;
signal FA3_l5_c43_S : std_logic;
signal FA3_l5_c43_Cout : std_logic;
signal FA4_l5_c43_S : std_logic;
signal FA4_l5_c43_Cout : std_logic;
signal FA1_l5_c44_S : std_logic;
signal FA1_l5_c44_Cout : std_logic;
signal FA2_l5_c44_S : std_logic;
signal FA2_l5_c44_Cout : std_logic;
signal FA3_l5_c44_S : std_logic;
signal FA3_l5_c44_Cout : std_logic;
signal HA1_l5_c44_S : std_logic;
signal HA1_l5_c44_Cout : std_logic;
signal FA1_l5_c45_S : std_logic;
signal FA1_l5_c45_Cout : std_logic;
signal FA2_l5_c45_S : std_logic;
signal FA2_l5_c45_Cout : std_logic;
signal FA3_l5_c45_S : std_logic;
signal FA3_l5_c45_Cout : std_logic;
signal FA1_l5_c46_S : std_logic;
signal FA1_l5_c46_Cout : std_logic;
signal FA2_l5_c46_S : std_logic;
signal FA2_l5_c46_Cout : std_logic;
signal HA1_l5_c46_S : std_logic;
signal HA1_l5_c46_Cout : std_logic;
signal FA1_l5_c47_S : std_logic;
signal FA1_l5_c47_Cout : std_logic;
signal FA2_l5_c47_S : std_logic;
signal FA2_l5_c47_Cout : std_logic;
signal FA1_l5_c48_S : std_logic;
signal FA1_l5_c48_Cout : std_logic;
signal HA1_l5_c48_S : std_logic;
signal HA1_l5_c48_Cout : std_logic;
signal FA1_l5_c49_S : std_logic;
signal FA1_l5_c49_Cout : std_logic;
signal HA1_l5_c50_S : std_logic;
signal HA1_l5_c50_Cout : std_logic;
signal HA1_l4_c10_S : std_logic;
signal HA1_l4_c10_Cout : std_logic;
signal HA1_l4_c11_S : std_logic;
signal HA1_l4_c11_Cout : std_logic;
signal FA1_l4_c12_S : std_logic;
signal FA1_l4_c12_Cout : std_logic;
signal HA1_l4_c12_S : std_logic;
signal HA1_l4_c12_Cout : std_logic;
signal FA1_l4_c13_S : std_logic;
signal FA1_l4_c13_Cout : std_logic;
signal HA1_l4_c13_S : std_logic;
signal HA1_l4_c13_Cout : std_logic;
signal FA1_l4_c14_S : std_logic;
signal FA1_l4_c14_Cout : std_logic;
signal FA2_l4_c14_S : std_logic;
signal FA2_l4_c14_Cout : std_logic;
signal HA1_l4_c14_S : std_logic;
signal HA1_l4_c14_Cout : std_logic;
signal FA1_l4_c15_S : std_logic;
signal FA1_l4_c15_Cout : std_logic;
signal FA2_l4_c15_S : std_logic;
signal FA2_l4_c15_Cout : std_logic;
signal HA1_l4_c15_S : std_logic;
signal HA1_l4_c15_Cout : std_logic;
signal FA1_l4_c16_S : std_logic;
signal FA1_l4_c16_Cout : std_logic;
signal FA2_l4_c16_S : std_logic;
signal FA2_l4_c16_Cout : std_logic;
signal FA3_l4_c16_S : std_logic;
signal FA3_l4_c16_Cout : std_logic;
signal FA1_l4_c17_S : std_logic;
signal FA1_l4_c17_Cout : std_logic;
signal FA2_l4_c17_S : std_logic;
signal FA2_l4_c17_Cout : std_logic;
signal FA3_l4_c17_S : std_logic;
signal FA3_l4_c17_Cout : std_logic;
signal FA1_l4_c18_S : std_logic;
signal FA1_l4_c18_Cout : std_logic;
signal FA2_l4_c18_S : std_logic;
signal FA2_l4_c18_Cout : std_logic;
signal FA3_l4_c18_S : std_logic;
signal FA3_l4_c18_Cout : std_logic;
signal FA1_l4_c19_S : std_logic;
signal FA1_l4_c19_Cout : std_logic;
signal FA2_l4_c19_S : std_logic;
signal FA2_l4_c19_Cout : std_logic;
signal FA3_l4_c19_S : std_logic;
signal FA3_l4_c19_Cout : std_logic;
signal FA1_l4_c20_S : std_logic;
signal FA1_l4_c20_Cout : std_logic;
signal FA2_l4_c20_S : std_logic;
signal FA2_l4_c20_Cout : std_logic;
signal FA3_l4_c20_S : std_logic;
signal FA3_l4_c20_Cout : std_logic;
signal FA1_l4_c21_S : std_logic;
signal FA1_l4_c21_Cout : std_logic;
signal FA2_l4_c21_S : std_logic;
signal FA2_l4_c21_Cout : std_logic;
signal FA3_l4_c21_S : std_logic;
signal FA3_l4_c21_Cout : std_logic;
signal FA1_l4_c22_S : std_logic;
signal FA1_l4_c22_Cout : std_logic;
signal FA2_l4_c22_S : std_logic;
signal FA2_l4_c22_Cout : std_logic;
signal FA3_l4_c22_S : std_logic;
signal FA3_l4_c22_Cout : std_logic;
signal FA1_l4_c23_S : std_logic;
signal FA1_l4_c23_Cout : std_logic;
signal FA2_l4_c23_S : std_logic;
signal FA2_l4_c23_Cout : std_logic;
signal FA3_l4_c23_S : std_logic;
signal FA3_l4_c23_Cout : std_logic;
signal FA1_l4_c24_S : std_logic;
signal FA1_l4_c24_Cout : std_logic;
signal FA2_l4_c24_S : std_logic;
signal FA2_l4_c24_Cout : std_logic;
signal FA3_l4_c24_S : std_logic;
signal FA3_l4_c24_Cout : std_logic;
signal FA1_l4_c25_S : std_logic;
signal FA1_l4_c25_Cout : std_logic;
signal FA2_l4_c25_S : std_logic;
signal FA2_l4_c25_Cout : std_logic;
signal FA3_l4_c25_S : std_logic;
signal FA3_l4_c25_Cout : std_logic;
signal FA1_l4_c26_S : std_logic;
signal FA1_l4_c26_Cout : std_logic;
signal FA2_l4_c26_S : std_logic;
signal FA2_l4_c26_Cout : std_logic;
signal FA3_l4_c26_S : std_logic;
signal FA3_l4_c26_Cout : std_logic;
signal FA1_l4_c27_S : std_logic;
signal FA1_l4_c27_Cout : std_logic;
signal FA2_l4_c27_S : std_logic;
signal FA2_l4_c27_Cout : std_logic;
signal FA3_l4_c27_S : std_logic;
signal FA3_l4_c27_Cout : std_logic;
signal FA1_l4_c28_S : std_logic;
signal FA1_l4_c28_Cout : std_logic;
signal FA2_l4_c28_S : std_logic;
signal FA2_l4_c28_Cout : std_logic;
signal FA3_l4_c28_S : std_logic;
signal FA3_l4_c28_Cout : std_logic;
signal FA1_l4_c29_S : std_logic;
signal FA1_l4_c29_Cout : std_logic;
signal FA2_l4_c29_S : std_logic;
signal FA2_l4_c29_Cout : std_logic;
signal FA3_l4_c29_S : std_logic;
signal FA3_l4_c29_Cout : std_logic;
signal FA1_l4_c30_S : std_logic;
signal FA1_l4_c30_Cout : std_logic;
signal FA2_l4_c30_S : std_logic;
signal FA2_l4_c30_Cout : std_logic;
signal FA3_l4_c30_S : std_logic;
signal FA3_l4_c30_Cout : std_logic;
signal FA1_l4_c31_S : std_logic;
signal FA1_l4_c31_Cout : std_logic;
signal FA2_l4_c31_S : std_logic;
signal FA2_l4_c31_Cout : std_logic;
signal FA3_l4_c31_S : std_logic;
signal FA3_l4_c31_Cout : std_logic;
signal FA1_l4_c32_S : std_logic;
signal FA1_l4_c32_Cout : std_logic;
signal FA2_l4_c32_S : std_logic;
signal FA2_l4_c32_Cout : std_logic;
signal FA3_l4_c32_S : std_logic;
signal FA3_l4_c32_Cout : std_logic;
signal FA1_l4_c33_S : std_logic;
signal FA1_l4_c33_Cout : std_logic;
signal FA2_l4_c33_S : std_logic;
signal FA2_l4_c33_Cout : std_logic;
signal FA3_l4_c33_S : std_logic;
signal FA3_l4_c33_Cout : std_logic;
signal FA1_l4_c34_S : std_logic;
signal FA1_l4_c34_Cout : std_logic;
signal FA2_l4_c34_S : std_logic;
signal FA2_l4_c34_Cout : std_logic;
signal FA3_l4_c34_S : std_logic;
signal FA3_l4_c34_Cout : std_logic;
signal FA1_l4_c35_S : std_logic;
signal FA1_l4_c35_Cout : std_logic;
signal FA2_l4_c35_S : std_logic;
signal FA2_l4_c35_Cout : std_logic;
signal FA3_l4_c35_S : std_logic;
signal FA3_l4_c35_Cout : std_logic;
signal FA1_l4_c36_S : std_logic;
signal FA1_l4_c36_Cout : std_logic;
signal FA2_l4_c36_S : std_logic;
signal FA2_l4_c36_Cout : std_logic;
signal FA3_l4_c36_S : std_logic;
signal FA3_l4_c36_Cout : std_logic;
signal FA1_l4_c37_S : std_logic;
signal FA1_l4_c37_Cout : std_logic;
signal FA2_l4_c37_S : std_logic;
signal FA2_l4_c37_Cout : std_logic;
signal FA3_l4_c37_S : std_logic;
signal FA3_l4_c37_Cout : std_logic;
signal FA1_l4_c38_S : std_logic;
signal FA1_l4_c38_Cout : std_logic;
signal FA2_l4_c38_S : std_logic;
signal FA2_l4_c38_Cout : std_logic;
signal FA3_l4_c38_S : std_logic;
signal FA3_l4_c38_Cout : std_logic;
signal FA1_l4_c39_S : std_logic;
signal FA1_l4_c39_Cout : std_logic;
signal FA2_l4_c39_S : std_logic;
signal FA2_l4_c39_Cout : std_logic;
signal FA3_l4_c39_S : std_logic;
signal FA3_l4_c39_Cout : std_logic;
signal FA1_l4_c40_S : std_logic;
signal FA1_l4_c40_Cout : std_logic;
signal FA2_l4_c40_S : std_logic;
signal FA2_l4_c40_Cout : std_logic;
signal FA3_l4_c40_S : std_logic;
signal FA3_l4_c40_Cout : std_logic;
signal FA1_l4_c41_S : std_logic;
signal FA1_l4_c41_Cout : std_logic;
signal FA2_l4_c41_S : std_logic;
signal FA2_l4_c41_Cout : std_logic;
signal FA3_l4_c41_S : std_logic;
signal FA3_l4_c41_Cout : std_logic;
signal FA1_l4_c42_S : std_logic;
signal FA1_l4_c42_Cout : std_logic;
signal FA2_l4_c42_S : std_logic;
signal FA2_l4_c42_Cout : std_logic;
signal FA3_l4_c42_S : std_logic;
signal FA3_l4_c42_Cout : std_logic;
signal FA1_l4_c43_S : std_logic;
signal FA1_l4_c43_Cout : std_logic;
signal FA2_l4_c43_S : std_logic;
signal FA2_l4_c43_Cout : std_logic;
signal FA3_l4_c43_S : std_logic;
signal FA3_l4_c43_Cout : std_logic;
signal FA1_l4_c44_S : std_logic;
signal FA1_l4_c44_Cout : std_logic;
signal FA2_l4_c44_S : std_logic;
signal FA2_l4_c44_Cout : std_logic;
signal FA3_l4_c44_S : std_logic;
signal FA3_l4_c44_Cout : std_logic;
signal FA1_l4_c45_S : std_logic;
signal FA1_l4_c45_Cout : std_logic;
signal FA2_l4_c45_S : std_logic;
signal FA2_l4_c45_Cout : std_logic;
signal FA3_l4_c45_S : std_logic;
signal FA3_l4_c45_Cout : std_logic;
signal FA1_l4_c46_S : std_logic;
signal FA1_l4_c46_Cout : std_logic;
signal FA2_l4_c46_S : std_logic;
signal FA2_l4_c46_Cout : std_logic;
signal FA3_l4_c46_S : std_logic;
signal FA3_l4_c46_Cout : std_logic;
signal FA1_l4_c47_S : std_logic;
signal FA1_l4_c47_Cout : std_logic;
signal FA2_l4_c47_S : std_logic;
signal FA2_l4_c47_Cout : std_logic;
signal FA3_l4_c47_S : std_logic;
signal FA3_l4_c47_Cout : std_logic;
signal FA1_l4_c48_S : std_logic;
signal FA1_l4_c48_Cout : std_logic;
signal FA2_l4_c48_S : std_logic;
signal FA2_l4_c48_Cout : std_logic;
signal FA3_l4_c48_S : std_logic;
signal FA3_l4_c48_Cout : std_logic;
signal FA1_l4_c49_S : std_logic;
signal FA1_l4_c49_Cout : std_logic;
signal FA2_l4_c49_S : std_logic;
signal FA2_l4_c49_Cout : std_logic;
signal FA3_l4_c49_S : std_logic;
signal FA3_l4_c49_Cout : std_logic;
signal FA1_l4_c50_S : std_logic;
signal FA1_l4_c50_Cout : std_logic;
signal FA2_l4_c50_S : std_logic;
signal FA2_l4_c50_Cout : std_logic;
signal FA3_l4_c50_S : std_logic;
signal FA3_l4_c50_Cout : std_logic;
signal FA1_l4_c51_S : std_logic;
signal FA1_l4_c51_Cout : std_logic;
signal FA2_l4_c51_S : std_logic;
signal FA2_l4_c51_Cout : std_logic;
signal FA3_l4_c51_S : std_logic;
signal FA3_l4_c51_Cout : std_logic;
signal FA1_l4_c52_S : std_logic;
signal FA1_l4_c52_Cout : std_logic;
signal FA2_l4_c52_S : std_logic;
signal FA2_l4_c52_Cout : std_logic;
signal HA1_l4_c52_S : std_logic;
signal HA1_l4_c52_Cout : std_logic;
signal FA1_l4_c53_S : std_logic;
signal FA1_l4_c53_Cout : std_logic;
signal FA2_l4_c53_S : std_logic;
signal FA2_l4_c53_Cout : std_logic;
signal FA1_l4_c54_S : std_logic;
signal FA1_l4_c54_Cout : std_logic;
signal HA1_l4_c54_S : std_logic;
signal HA1_l4_c54_Cout : std_logic;
signal FA1_l4_c55_S : std_logic;
signal FA1_l4_c55_Cout : std_logic;
signal HA1_l4_c56_S : std_logic;
signal HA1_l4_c56_Cout : std_logic;
signal HA1_l3_c6_S : std_logic;
signal HA1_l3_c6_Cout : std_logic;
signal HA1_l3_c7_S : std_logic;
signal HA1_l3_c7_Cout : std_logic;
signal FA1_l3_c8_S : std_logic;
signal FA1_l3_c8_Cout : std_logic;
signal HA1_l3_c8_S : std_logic;
signal HA1_l3_c8_Cout : std_logic;
signal FA1_l3_c9_S : std_logic;
signal FA1_l3_c9_Cout : std_logic;
signal HA1_l3_c9_S : std_logic;
signal HA1_l3_c9_Cout : std_logic;
signal FA1_l3_c10_S : std_logic;
signal FA1_l3_c10_Cout : std_logic;
signal FA2_l3_c10_S : std_logic;
signal FA2_l3_c10_Cout : std_logic;
signal FA1_l3_c11_S : std_logic;
signal FA1_l3_c11_Cout : std_logic;
signal FA2_l3_c11_S : std_logic;
signal FA2_l3_c11_Cout : std_logic;
signal FA1_l3_c12_S : std_logic;
signal FA1_l3_c12_Cout : std_logic;
signal FA2_l3_c12_S : std_logic;
signal FA2_l3_c12_Cout : std_logic;
signal FA1_l3_c13_S : std_logic;
signal FA1_l3_c13_Cout : std_logic;
signal FA2_l3_c13_S : std_logic;
signal FA2_l3_c13_Cout : std_logic;
signal FA1_l3_c14_S : std_logic;
signal FA1_l3_c14_Cout : std_logic;
signal FA2_l3_c14_S : std_logic;
signal FA2_l3_c14_Cout : std_logic;
signal FA1_l3_c15_S : std_logic;
signal FA1_l3_c15_Cout : std_logic;
signal FA2_l3_c15_S : std_logic;
signal FA2_l3_c15_Cout : std_logic;
signal FA1_l3_c16_S : std_logic;
signal FA1_l3_c16_Cout : std_logic;
signal FA2_l3_c16_S : std_logic;
signal FA2_l3_c16_Cout : std_logic;
signal FA1_l3_c17_S : std_logic;
signal FA1_l3_c17_Cout : std_logic;
signal FA2_l3_c17_S : std_logic;
signal FA2_l3_c17_Cout : std_logic;
signal FA1_l3_c18_S : std_logic;
signal FA1_l3_c18_Cout : std_logic;
signal FA2_l3_c18_S : std_logic;
signal FA2_l3_c18_Cout : std_logic;
signal FA1_l3_c19_S : std_logic;
signal FA1_l3_c19_Cout : std_logic;
signal FA2_l3_c19_S : std_logic;
signal FA2_l3_c19_Cout : std_logic;
signal FA1_l3_c20_S : std_logic;
signal FA1_l3_c20_Cout : std_logic;
signal FA2_l3_c20_S : std_logic;
signal FA2_l3_c20_Cout : std_logic;
signal FA1_l3_c21_S : std_logic;
signal FA1_l3_c21_Cout : std_logic;
signal FA2_l3_c21_S : std_logic;
signal FA2_l3_c21_Cout : std_logic;
signal FA1_l3_c22_S : std_logic;
signal FA1_l3_c22_Cout : std_logic;
signal FA2_l3_c22_S : std_logic;
signal FA2_l3_c22_Cout : std_logic;
signal FA1_l3_c23_S : std_logic;
signal FA1_l3_c23_Cout : std_logic;
signal FA2_l3_c23_S : std_logic;
signal FA2_l3_c23_Cout : std_logic;
signal FA1_l3_c24_S : std_logic;
signal FA1_l3_c24_Cout : std_logic;
signal FA2_l3_c24_S : std_logic;
signal FA2_l3_c24_Cout : std_logic;
signal FA1_l3_c25_S : std_logic;
signal FA1_l3_c25_Cout : std_logic;
signal FA2_l3_c25_S : std_logic;
signal FA2_l3_c25_Cout : std_logic;
signal FA1_l3_c26_S : std_logic;
signal FA1_l3_c26_Cout : std_logic;
signal FA2_l3_c26_S : std_logic;
signal FA2_l3_c26_Cout : std_logic;
signal FA1_l3_c27_S : std_logic;
signal FA1_l3_c27_Cout : std_logic;
signal FA2_l3_c27_S : std_logic;
signal FA2_l3_c27_Cout : std_logic;
signal FA1_l3_c28_S : std_logic;
signal FA1_l3_c28_Cout : std_logic;
signal FA2_l3_c28_S : std_logic;
signal FA2_l3_c28_Cout : std_logic;
signal FA1_l3_c29_S : std_logic;
signal FA1_l3_c29_Cout : std_logic;
signal FA2_l3_c29_S : std_logic;
signal FA2_l3_c29_Cout : std_logic;
signal FA1_l3_c30_S : std_logic;
signal FA1_l3_c30_Cout : std_logic;
signal FA2_l3_c30_S : std_logic;
signal FA2_l3_c30_Cout : std_logic;
signal FA1_l3_c31_S : std_logic;
signal FA1_l3_c31_Cout : std_logic;
signal FA2_l3_c31_S : std_logic;
signal FA2_l3_c31_Cout : std_logic;
signal FA1_l3_c32_S : std_logic;
signal FA1_l3_c32_Cout : std_logic;
signal FA2_l3_c32_S : std_logic;
signal FA2_l3_c32_Cout : std_logic;
signal FA1_l3_c33_S : std_logic;
signal FA1_l3_c33_Cout : std_logic;
signal FA2_l3_c33_S : std_logic;
signal FA2_l3_c33_Cout : std_logic;
signal FA1_l3_c34_S : std_logic;
signal FA1_l3_c34_Cout : std_logic;
signal FA2_l3_c34_S : std_logic;
signal FA2_l3_c34_Cout : std_logic;
signal FA1_l3_c35_S : std_logic;
signal FA1_l3_c35_Cout : std_logic;
signal FA2_l3_c35_S : std_logic;
signal FA2_l3_c35_Cout : std_logic;
signal FA1_l3_c36_S : std_logic;
signal FA1_l3_c36_Cout : std_logic;
signal FA2_l3_c36_S : std_logic;
signal FA2_l3_c36_Cout : std_logic;
signal FA1_l3_c37_S : std_logic;
signal FA1_l3_c37_Cout : std_logic;
signal FA2_l3_c37_S : std_logic;
signal FA2_l3_c37_Cout : std_logic;
signal FA1_l3_c38_S : std_logic;
signal FA1_l3_c38_Cout : std_logic;
signal FA2_l3_c38_S : std_logic;
signal FA2_l3_c38_Cout : std_logic;
signal FA1_l3_c39_S : std_logic;
signal FA1_l3_c39_Cout : std_logic;
signal FA2_l3_c39_S : std_logic;
signal FA2_l3_c39_Cout : std_logic;
signal FA1_l3_c40_S : std_logic;
signal FA1_l3_c40_Cout : std_logic;
signal FA2_l3_c40_S : std_logic;
signal FA2_l3_c40_Cout : std_logic;
signal FA1_l3_c41_S : std_logic;
signal FA1_l3_c41_Cout : std_logic;
signal FA2_l3_c41_S : std_logic;
signal FA2_l3_c41_Cout : std_logic;
signal FA1_l3_c42_S : std_logic;
signal FA1_l3_c42_Cout : std_logic;
signal FA2_l3_c42_S : std_logic;
signal FA2_l3_c42_Cout : std_logic;
signal FA1_l3_c43_S : std_logic;
signal FA1_l3_c43_Cout : std_logic;
signal FA2_l3_c43_S : std_logic;
signal FA2_l3_c43_Cout : std_logic;
signal FA1_l3_c44_S : std_logic;
signal FA1_l3_c44_Cout : std_logic;
signal FA2_l3_c44_S : std_logic;
signal FA2_l3_c44_Cout : std_logic;
signal FA1_l3_c45_S : std_logic;
signal FA1_l3_c45_Cout : std_logic;
signal FA2_l3_c45_S : std_logic;
signal FA2_l3_c45_Cout : std_logic;
signal FA1_l3_c46_S : std_logic;
signal FA1_l3_c46_Cout : std_logic;
signal FA2_l3_c46_S : std_logic;
signal FA2_l3_c46_Cout : std_logic;
signal FA1_l3_c47_S : std_logic;
signal FA1_l3_c47_Cout : std_logic;
signal FA2_l3_c47_S : std_logic;
signal FA2_l3_c47_Cout : std_logic;
signal FA1_l3_c48_S : std_logic;
signal FA1_l3_c48_Cout : std_logic;
signal FA2_l3_c48_S : std_logic;
signal FA2_l3_c48_Cout : std_logic;
signal FA1_l3_c49_S : std_logic;
signal FA1_l3_c49_Cout : std_logic;
signal FA2_l3_c49_S : std_logic;
signal FA2_l3_c49_Cout : std_logic;
signal FA1_l3_c50_S : std_logic;
signal FA1_l3_c50_Cout : std_logic;
signal FA2_l3_c50_S : std_logic;
signal FA2_l3_c50_Cout : std_logic;
signal FA1_l3_c51_S : std_logic;
signal FA1_l3_c51_Cout : std_logic;
signal FA2_l3_c51_S : std_logic;
signal FA2_l3_c51_Cout : std_logic;
signal FA1_l3_c52_S : std_logic;
signal FA1_l3_c52_Cout : std_logic;
signal FA2_l3_c52_S : std_logic;
signal FA2_l3_c52_Cout : std_logic;
signal FA1_l3_c53_S : std_logic;
signal FA1_l3_c53_Cout : std_logic;
signal FA2_l3_c53_S : std_logic;
signal FA2_l3_c53_Cout : std_logic;
signal FA1_l3_c54_S : std_logic;
signal FA1_l3_c54_Cout : std_logic;
signal FA2_l3_c54_S : std_logic;
signal FA2_l3_c54_Cout : std_logic;
signal FA1_l3_c55_S : std_logic;
signal FA1_l3_c55_Cout : std_logic;
signal FA2_l3_c55_S : std_logic;
signal FA2_l3_c55_Cout : std_logic;
signal FA1_l3_c56_S : std_logic;
signal FA1_l3_c56_Cout : std_logic;
signal FA2_l3_c56_S : std_logic;
signal FA2_l3_c56_Cout : std_logic;
signal FA1_l3_c57_S : std_logic;
signal FA1_l3_c57_Cout : std_logic;
signal FA2_l3_c57_S : std_logic;
signal FA2_l3_c57_Cout : std_logic;
signal FA1_l3_c58_S : std_logic;
signal FA1_l3_c58_Cout : std_logic;
signal HA1_l3_c58_S : std_logic;
signal HA1_l3_c58_Cout : std_logic;
signal FA1_l3_c59_S : std_logic;
signal FA1_l3_c59_Cout : std_logic;
signal HA1_l3_c60_S : std_logic;
signal HA1_l3_c60_Cout : std_logic;
signal HA1_l2_c4_S : std_logic;
signal HA1_l2_c4_Cout : std_logic;
signal HA1_l2_c5_S : std_logic;
signal HA1_l2_c5_Cout : std_logic;
signal FA1_l2_c6_S : std_logic;
signal FA1_l2_c6_Cout : std_logic;
signal FA1_l2_c7_S : std_logic;
signal FA1_l2_c7_Cout : std_logic;
signal FA1_l2_c8_S : std_logic;
signal FA1_l2_c8_Cout : std_logic;
signal FA1_l2_c9_S : std_logic;
signal FA1_l2_c9_Cout : std_logic;
signal FA1_l2_c10_S : std_logic;
signal FA1_l2_c10_Cout : std_logic;
signal FA1_l2_c11_S : std_logic;
signal FA1_l2_c11_Cout : std_logic;
signal FA1_l2_c12_S : std_logic;
signal FA1_l2_c12_Cout : std_logic;
signal FA1_l2_c13_S : std_logic;
signal FA1_l2_c13_Cout : std_logic;
signal FA1_l2_c14_S : std_logic;
signal FA1_l2_c14_Cout : std_logic;
signal FA1_l2_c15_S : std_logic;
signal FA1_l2_c15_Cout : std_logic;
signal FA1_l2_c16_S : std_logic;
signal FA1_l2_c16_Cout : std_logic;
signal FA1_l2_c17_S : std_logic;
signal FA1_l2_c17_Cout : std_logic;
signal FA1_l2_c18_S : std_logic;
signal FA1_l2_c18_Cout : std_logic;
signal FA1_l2_c19_S : std_logic;
signal FA1_l2_c19_Cout : std_logic;
signal FA1_l2_c20_S : std_logic;
signal FA1_l2_c20_Cout : std_logic;
signal FA1_l2_c21_S : std_logic;
signal FA1_l2_c21_Cout : std_logic;
signal FA1_l2_c22_S : std_logic;
signal FA1_l2_c22_Cout : std_logic;
signal FA1_l2_c23_S : std_logic;
signal FA1_l2_c23_Cout : std_logic;
signal FA1_l2_c24_S : std_logic;
signal FA1_l2_c24_Cout : std_logic;
signal FA1_l2_c25_S : std_logic;
signal FA1_l2_c25_Cout : std_logic;
signal FA1_l2_c26_S : std_logic;
signal FA1_l2_c26_Cout : std_logic;
signal FA1_l2_c27_S : std_logic;
signal FA1_l2_c27_Cout : std_logic;
signal FA1_l2_c28_S : std_logic;
signal FA1_l2_c28_Cout : std_logic;
signal FA1_l2_c29_S : std_logic;
signal FA1_l2_c29_Cout : std_logic;
signal FA1_l2_c30_S : std_logic;
signal FA1_l2_c30_Cout : std_logic;
signal FA1_l2_c31_S : std_logic;
signal FA1_l2_c31_Cout : std_logic;
signal FA1_l2_c32_S : std_logic;
signal FA1_l2_c32_Cout : std_logic;
signal FA1_l2_c33_S : std_logic;
signal FA1_l2_c33_Cout : std_logic;
signal FA1_l2_c34_S : std_logic;
signal FA1_l2_c34_Cout : std_logic;
signal FA1_l2_c35_S : std_logic;
signal FA1_l2_c35_Cout : std_logic;
signal FA1_l2_c36_S : std_logic;
signal FA1_l2_c36_Cout : std_logic;
signal FA1_l2_c37_S : std_logic;
signal FA1_l2_c37_Cout : std_logic;
signal FA1_l2_c38_S : std_logic;
signal FA1_l2_c38_Cout : std_logic;
signal FA1_l2_c39_S : std_logic;
signal FA1_l2_c39_Cout : std_logic;
signal FA1_l2_c40_S : std_logic;
signal FA1_l2_c40_Cout : std_logic;
signal FA1_l2_c41_S : std_logic;
signal FA1_l2_c41_Cout : std_logic;
signal FA1_l2_c42_S : std_logic;
signal FA1_l2_c42_Cout : std_logic;
signal FA1_l2_c43_S : std_logic;
signal FA1_l2_c43_Cout : std_logic;
signal FA1_l2_c44_S : std_logic;
signal FA1_l2_c44_Cout : std_logic;
signal FA1_l2_c45_S : std_logic;
signal FA1_l2_c45_Cout : std_logic;
signal FA1_l2_c46_S : std_logic;
signal FA1_l2_c46_Cout : std_logic;
signal FA1_l2_c47_S : std_logic;
signal FA1_l2_c47_Cout : std_logic;
signal FA1_l2_c48_S : std_logic;
signal FA1_l2_c48_Cout : std_logic;
signal FA1_l2_c49_S : std_logic;
signal FA1_l2_c49_Cout : std_logic;
signal FA1_l2_c50_S : std_logic;
signal FA1_l2_c50_Cout : std_logic;
signal FA1_l2_c51_S : std_logic;
signal FA1_l2_c51_Cout : std_logic;
signal FA1_l2_c52_S : std_logic;
signal FA1_l2_c52_Cout : std_logic;
signal FA1_l2_c53_S : std_logic;
signal FA1_l2_c53_Cout : std_logic;
signal FA1_l2_c54_S : std_logic;
signal FA1_l2_c54_Cout : std_logic;
signal FA1_l2_c55_S : std_logic;
signal FA1_l2_c55_Cout : std_logic;
signal FA1_l2_c56_S : std_logic;
signal FA1_l2_c56_Cout : std_logic;
signal FA1_l2_c57_S : std_logic;
signal FA1_l2_c57_Cout : std_logic;
signal FA1_l2_c58_S : std_logic;
signal FA1_l2_c58_Cout : std_logic;
signal FA1_l2_c59_S : std_logic;
signal FA1_l2_c59_Cout : std_logic;
signal FA1_l2_c60_S : std_logic;
signal FA1_l2_c60_Cout : std_logic;
signal FA1_l2_c61_S : std_logic;
signal FA1_l2_c61_Cout : std_logic;
signal HA1_l2_c62_S : std_logic;
signal HA1_l2_c62_Cout : std_logic;
signal HA1_l1_c2_S : std_logic;
signal HA1_l1_c2_Cout : std_logic;
signal HA1_l1_c3_S : std_logic;
signal HA1_l1_c3_Cout : std_logic;
signal FA1_l1_c4_S : std_logic;
signal FA1_l1_c4_Cout : std_logic;
signal FA1_l1_c5_S : std_logic;
signal FA1_l1_c5_Cout : std_logic;
signal FA1_l1_c6_S : std_logic;
signal FA1_l1_c6_Cout : std_logic;
signal FA1_l1_c7_S : std_logic;
signal FA1_l1_c7_Cout : std_logic;
signal FA1_l1_c8_S : std_logic;
signal FA1_l1_c8_Cout : std_logic;
signal FA1_l1_c9_S : std_logic;
signal FA1_l1_c9_Cout : std_logic;
signal FA1_l1_c10_S : std_logic;
signal FA1_l1_c10_Cout : std_logic;
signal FA1_l1_c11_S : std_logic;
signal FA1_l1_c11_Cout : std_logic;
signal FA1_l1_c12_S : std_logic;
signal FA1_l1_c12_Cout : std_logic;
signal FA1_l1_c13_S : std_logic;
signal FA1_l1_c13_Cout : std_logic;
signal FA1_l1_c14_S : std_logic;
signal FA1_l1_c14_Cout : std_logic;
signal FA1_l1_c15_S : std_logic;
signal FA1_l1_c15_Cout : std_logic;
signal FA1_l1_c16_S : std_logic;
signal FA1_l1_c16_Cout : std_logic;
signal FA1_l1_c17_S : std_logic;
signal FA1_l1_c17_Cout : std_logic;
signal FA1_l1_c18_S : std_logic;
signal FA1_l1_c18_Cout : std_logic;
signal FA1_l1_c19_S : std_logic;
signal FA1_l1_c19_Cout : std_logic;
signal FA1_l1_c20_S : std_logic;
signal FA1_l1_c20_Cout : std_logic;
signal FA1_l1_c21_S : std_logic;
signal FA1_l1_c21_Cout : std_logic;
signal FA1_l1_c22_S : std_logic;
signal FA1_l1_c22_Cout : std_logic;
signal FA1_l1_c23_S : std_logic;
signal FA1_l1_c23_Cout : std_logic;
signal FA1_l1_c24_S : std_logic;
signal FA1_l1_c24_Cout : std_logic;
signal FA1_l1_c25_S : std_logic;
signal FA1_l1_c25_Cout : std_logic;
signal FA1_l1_c26_S : std_logic;
signal FA1_l1_c26_Cout : std_logic;
signal FA1_l1_c27_S : std_logic;
signal FA1_l1_c27_Cout : std_logic;
signal FA1_l1_c28_S : std_logic;
signal FA1_l1_c28_Cout : std_logic;
signal FA1_l1_c29_S : std_logic;
signal FA1_l1_c29_Cout : std_logic;
signal FA1_l1_c30_S : std_logic;
signal FA1_l1_c30_Cout : std_logic;
signal FA1_l1_c31_S : std_logic;
signal FA1_l1_c31_Cout : std_logic;
signal FA1_l1_c32_S : std_logic;
signal FA1_l1_c32_Cout : std_logic;
signal FA1_l1_c33_S : std_logic;
signal FA1_l1_c33_Cout : std_logic;
signal FA1_l1_c34_S : std_logic;
signal FA1_l1_c34_Cout : std_logic;
signal FA1_l1_c35_S : std_logic;
signal FA1_l1_c35_Cout : std_logic;
signal FA1_l1_c36_S : std_logic;
signal FA1_l1_c36_Cout : std_logic;
signal FA1_l1_c37_S : std_logic;
signal FA1_l1_c37_Cout : std_logic;
signal FA1_l1_c38_S : std_logic;
signal FA1_l1_c38_Cout : std_logic;
signal FA1_l1_c39_S : std_logic;
signal FA1_l1_c39_Cout : std_logic;
signal FA1_l1_c40_S : std_logic;
signal FA1_l1_c40_Cout : std_logic;
signal FA1_l1_c41_S : std_logic;
signal FA1_l1_c41_Cout : std_logic;
signal FA1_l1_c42_S : std_logic;
signal FA1_l1_c42_Cout : std_logic;
signal FA1_l1_c43_S : std_logic;
signal FA1_l1_c43_Cout : std_logic;
signal FA1_l1_c44_S : std_logic;
signal FA1_l1_c44_Cout : std_logic;
signal FA1_l1_c45_S : std_logic;
signal FA1_l1_c45_Cout : std_logic;
signal FA1_l1_c46_S : std_logic;
signal FA1_l1_c46_Cout : std_logic;
signal FA1_l1_c47_S : std_logic;
signal FA1_l1_c47_Cout : std_logic;
signal FA1_l1_c48_S : std_logic;
signal FA1_l1_c48_Cout : std_logic;
signal FA1_l1_c49_S : std_logic;
signal FA1_l1_c49_Cout : std_logic;
signal FA1_l1_c50_S : std_logic;
signal FA1_l1_c50_Cout : std_logic;
signal FA1_l1_c51_S : std_logic;
signal FA1_l1_c51_Cout : std_logic;
signal FA1_l1_c52_S : std_logic;
signal FA1_l1_c52_Cout : std_logic;
signal FA1_l1_c53_S : std_logic;
signal FA1_l1_c53_Cout : std_logic;
signal FA1_l1_c54_S : std_logic;
signal FA1_l1_c54_Cout : std_logic;
signal FA1_l1_c55_S : std_logic;
signal FA1_l1_c55_Cout : std_logic;
signal FA1_l1_c56_S : std_logic;
signal FA1_l1_c56_Cout : std_logic;
signal FA1_l1_c57_S : std_logic;
signal FA1_l1_c57_Cout : std_logic;
signal FA1_l1_c58_S : std_logic;
signal FA1_l1_c58_Cout : std_logic;
signal FA1_l1_c59_S : std_logic;
signal FA1_l1_c59_Cout : std_logic;
signal FA1_l1_c60_S : std_logic;
signal FA1_l1_c60_Cout : std_logic;
signal FA1_l1_c61_S : std_logic;
signal FA1_l1_c61_Cout : std_logic;
signal FA1_l1_c62_S : std_logic;
signal FA1_l1_c62_Cout : std_logic;
signal FA1_l1_c63_S : std_logic;
signal FA1_l1_c63_Cout : std_logic;	

signal sum_1 : std_logic_vector(63 downto 0);
signal sum_2 : std_logic_vector(63 downto 0);

signal sum : std_logic_vector(63 downto 0);

begin

	PP0_neg <= NOT PP0(32);
	PP1_neg <= NOT PP1(32);
	PP2_neg <= NOT PP2(32);
	PP3_neg <= NOT PP3(32);
	PP4_neg <= NOT PP4(32);
	PP5_neg <= NOT PP5(32);
	PP6_neg <= NOT PP6(32);
	PP7_neg <= NOT PP7(32);
	PP8_neg <= NOT PP8(32);
	PP9_neg <= NOT PP9(32);
	PP10_neg <= NOT PP10(32);
	PP11_neg <= NOT PP11(32);
	PP12_neg <= NOT PP12(32);
	PP13_neg <= NOT PP13(32);
	PP14_neg <= NOT PP14(32);
	PP15_neg <= NOT PP15(32);

	sum_1(1 DOWNTO 0) <= PP0(1 DOWNTO 0);
	sum_1(2) <= HA1_l1_c2_S;
	sum_1(3) <= HA1_l1_c3_S;
	sum_1(4) <= FA1_l1_c4_S;
	sum_1(5) <= FA1_l1_c5_S;
	sum_1(6) <= FA1_l1_c6_S;
	sum_1(7) <= FA1_l1_c7_S;
	sum_1(8) <= FA1_l1_c8_S;
	sum_1(9) <= FA1_l1_c9_S;
	sum_1(10) <= FA1_l1_c10_S;
	sum_1(11) <= FA1_l1_c11_S;
	sum_1(12) <= FA1_l1_c12_S;
	sum_1(13) <= FA1_l1_c13_S;
	sum_1(14) <= FA1_l1_c14_S;
	sum_1(15) <= FA1_l1_c15_S;
	sum_1(16) <= FA1_l1_c16_S;
	sum_1(17) <= FA1_l1_c17_S;
	sum_1(18) <= FA1_l1_c18_S;
	sum_1(19) <= FA1_l1_c19_S;
	sum_1(20) <= FA1_l1_c20_S;
	sum_1(21) <= FA1_l1_c21_S;
	sum_1(22) <= FA1_l1_c22_S;
	sum_1(23) <= FA1_l1_c23_S;
	sum_1(24) <= FA1_l1_c24_S;
	sum_1(25) <= FA1_l1_c25_S;
	sum_1(26) <= FA1_l1_c26_S;
	sum_1(27) <= FA1_l1_c27_S;
	sum_1(28) <= FA1_l1_c28_S;
	sum_1(29) <= FA1_l1_c29_S;
	sum_1(30) <= FA1_l1_c30_S;
	sum_1(31) <= FA1_l1_c31_S;
	sum_1(32) <= FA1_l1_c32_S;
	sum_1(33) <= FA1_l1_c33_S;
	sum_1(34) <= FA1_l1_c34_S;
	sum_1(35) <= FA1_l1_c35_S;
	sum_1(36) <= FA1_l1_c36_S;
	sum_1(37) <= FA1_l1_c37_S;
	sum_1(38) <= FA1_l1_c38_S;
	sum_1(39) <= FA1_l1_c39_S;
	sum_1(40) <= FA1_l1_c40_S;
	sum_1(41) <= FA1_l1_c41_S;
	sum_1(42) <= FA1_l1_c42_S;
	sum_1(43) <= FA1_l1_c43_S;
	sum_1(44) <= FA1_l1_c44_S;
	sum_1(45) <= FA1_l1_c45_S;
	sum_1(46) <= FA1_l1_c46_S;
	sum_1(47) <= FA1_l1_c47_S;
	sum_1(48) <= FA1_l1_c48_S;
	sum_1(49) <= FA1_l1_c49_S;
	sum_1(50) <= FA1_l1_c50_S;
	sum_1(51) <= FA1_l1_c51_S;
	sum_1(52) <= FA1_l1_c52_S;
	sum_1(53) <= FA1_l1_c53_S;
	sum_1(54) <= FA1_l1_c54_S;
	sum_1(55) <= FA1_l1_c55_S;
	sum_1(56) <= FA1_l1_c56_S;
	sum_1(57) <= FA1_l1_c57_S;
	sum_1(58) <= FA1_l1_c58_S;
	sum_1(59) <= FA1_l1_c59_S;
	sum_1(60) <= FA1_l1_c60_S;
	sum_1(61) <= FA1_l1_c61_S;
	sum_1(62) <= FA1_l1_c62_S;
	sum_1(63) <= FA1_l1_c63_S;

	sum_2(0) <= PP0(32);
	sum_2(1) <= '0';
	sum_2(2) <= PP1(32);
	sum_2(3) <= HA1_l1_c2_Cout;
	sum_2(4) <= HA1_l1_c3_Cout;
	sum_2(5) <= FA1_l1_c4_Cout;
	sum_2(6) <= FA1_l1_c5_Cout;
	sum_2(7) <= FA1_l1_c6_Cout;
	sum_2(8) <= FA1_l1_c7_Cout;
	sum_2(9) <= FA1_l1_c8_Cout;
	sum_2(10) <= FA1_l1_c9_Cout;
	sum_2(11) <= FA1_l1_c10_Cout;
	sum_2(12) <= FA1_l1_c11_Cout;
	sum_2(13) <= FA1_l1_c12_Cout;
	sum_2(14) <= FA1_l1_c13_Cout;
	sum_2(15) <= FA1_l1_c14_Cout;
	sum_2(16) <= FA1_l1_c15_Cout;
	sum_2(17) <= FA1_l1_c16_Cout;
	sum_2(18) <= FA1_l1_c17_Cout;
	sum_2(19) <= FA1_l1_c18_Cout;
	sum_2(20) <= FA1_l1_c19_Cout;
	sum_2(21) <= FA1_l1_c20_Cout;
	sum_2(22) <= FA1_l1_c21_Cout;
	sum_2(23) <= FA1_l1_c22_Cout;
	sum_2(24) <= FA1_l1_c23_Cout;
	sum_2(25) <= FA1_l1_c24_Cout;
	sum_2(26) <= FA1_l1_c25_Cout;
	sum_2(27) <= FA1_l1_c26_Cout;
	sum_2(28) <= FA1_l1_c27_Cout;
	sum_2(29) <= FA1_l1_c28_Cout;
	sum_2(30) <= FA1_l1_c29_Cout;
	sum_2(31) <= FA1_l1_c30_Cout;
	sum_2(32) <= FA1_l1_c31_Cout;
	sum_2(33) <= FA1_l1_c32_Cout;
	sum_2(34) <= FA1_l1_c33_Cout;
	sum_2(35) <= FA1_l1_c34_Cout;
	sum_2(36) <= FA1_l1_c35_Cout;
	sum_2(37) <= FA1_l1_c36_Cout;
	sum_2(38) <= FA1_l1_c37_Cout;
	sum_2(39) <= FA1_l1_c38_Cout;
	sum_2(40) <= FA1_l1_c39_Cout;
	sum_2(41) <= FA1_l1_c40_Cout;
	sum_2(42) <= FA1_l1_c41_Cout;
	sum_2(43) <= FA1_l1_c42_Cout;
	sum_2(44) <= FA1_l1_c43_Cout;
	sum_2(45) <= FA1_l1_c44_Cout;
	sum_2(46) <= FA1_l1_c45_Cout;
	sum_2(47) <= FA1_l1_c46_Cout;
	sum_2(48) <= FA1_l1_c47_Cout;
	sum_2(49) <= FA1_l1_c48_Cout;
	sum_2(50) <= FA1_l1_c49_Cout;
	sum_2(51) <= FA1_l1_c50_Cout;
	sum_2(52) <= FA1_l1_c51_Cout;
	sum_2(53) <= FA1_l1_c52_Cout;
	sum_2(54) <= FA1_l1_c53_Cout;
	sum_2(55) <= FA1_l1_c54_Cout;
	sum_2(56) <= FA1_l1_c55_Cout;
	sum_2(57) <= FA1_l1_c56_Cout;
	sum_2(58) <= FA1_l1_c57_Cout;
	sum_2(59) <= FA1_l1_c58_Cout;
	sum_2(60) <= FA1_l1_c59_Cout;
	sum_2(61) <= FA1_l1_c60_Cout;
	sum_2(62) <= FA1_l1_c61_Cout;
	sum_2(63) <= FA1_l1_c62_Cout;

	partial_product_generator  : PP_gen 
	PORT MAP ( A => A,
				  B => B, 
				  PP0	=> PP0, 
				  PP1	=> PP1, 
				  PP2	=> PP2, 
				  PP3	=> PP3, 
				  PP4	=> PP4, 
				  PP5	=> PP5, 
				  PP6	=> PP6, 
				  PP7	=> PP7, 
				  PP8	=> PP8, 
				  PP9	=> PP9,
				  PP10 => PP10, 
				  PP11 => PP11, 
				  PP12 => PP12,
				  PP13 => PP13,
				  PP14 => PP14, 
				  PP15 => PP15, 
				  PP16 => PP16);

	HA1_l6_c24  : HA 
	PORT MAP ( A =>	PP0(24), B =>	PP1(22), S =>	HA1_l6_c24_S, COUT 	=>	HA1_l6_c24_Cout );

	HA1_l6_c25  : HA 
	PORT MAP ( A =>	PP0(25), B =>	PP1(23), S =>	HA1_l6_c25_S, COUT 	=>	HA1_l6_c25_Cout );

	FA1_l6_c26  : FA 
	PORT MAP ( A =>	PP0(26), B =>	PP1(24), CIN 	=>	PP2(22), S =>	FA1_l6_c26_S, COUT 	=>	FA1_l6_c26_Cout );

	HA1_l6_c26  : HA 
	PORT MAP ( A =>	PP3(20), B =>	PP4(18), S =>	HA1_l6_c26_S, COUT 	=>	HA1_l6_c26_Cout );

	FA1_l6_c27  : FA 
	PORT MAP ( A =>	PP0(27), B =>	PP1(25), CIN 	=>	PP2(23), S =>	FA1_l6_c27_S, COUT 	=>	FA1_l6_c27_Cout );

	HA1_l6_c27  : HA 
	PORT MAP ( A =>	PP3(21), B =>	PP4(19), S =>	HA1_l6_c27_S, COUT 	=>	HA1_l6_c27_Cout );

	FA1_l6_c28  : FA 
	PORT MAP ( A =>	PP0(28), B =>	PP1(26), CIN 	=>	PP2(24), S =>	FA1_l6_c28_S, COUT 	=>	FA1_l6_c28_Cout );

	FA2_l6_c28  : FA 
	PORT MAP ( A =>	PP3(22), B =>	PP4(20), CIN 	=>	PP5(18), S =>	FA2_l6_c28_S, COUT 	=>	FA2_l6_c28_Cout );

	HA1_l6_c28  : HA 
	PORT MAP ( A =>	PP6(16), B =>	PP7(14), S =>	HA1_l6_c28_S, COUT 	=>	HA1_l6_c28_Cout );

	FA1_l6_c29  : FA 
	PORT MAP ( A =>	PP0(29), B =>	PP1(27), CIN 	=>	PP2(25), S =>	FA1_l6_c29_S, COUT 	=>	FA1_l6_c29_Cout );

	FA2_l6_c29  : FA 
	PORT MAP ( A =>	PP3(23), B =>	PP4(21), CIN 	=>	PP5(19), S =>	FA2_l6_c29_S, COUT 	=>	FA2_l6_c29_Cout );

	HA1_l6_c29  : HA 
	PORT MAP ( A =>	PP6(17), B =>	PP7(15), S =>	HA1_l6_c29_S, COUT 	=>	HA1_l6_c29_Cout );

	FA1_l6_c30  : FA 
	PORT MAP ( A =>	PP0(30), B =>	PP1(28), CIN 	=>	PP2(26), S =>	FA1_l6_c30_S, COUT 	=>	FA1_l6_c30_Cout );

	FA2_l6_c30  : FA 
	PORT MAP ( A =>	PP3(24), B =>	PP4(22), CIN 	=>	PP5(20), S =>	FA2_l6_c30_S, COUT 	=>	FA2_l6_c30_Cout );

	FA3_l6_c30  : FA 
	PORT MAP ( A =>	PP6(18), B =>	PP7(16), CIN 	=>	PP8(14), S =>	FA3_l6_c30_S, COUT 	=>	FA3_l6_c30_Cout );

	HA1_l6_c30  : HA 
	PORT MAP ( A =>	PP9(12), B =>	PP10(10), S =>	HA1_l6_c30_S, COUT 	=>	HA1_l6_c30_Cout );

	FA1_l6_c31  : FA 
	PORT MAP ( A =>	PP0(31), B =>	PP1(29), CIN 	=>	PP2(27), S =>	FA1_l6_c31_S, COUT 	=>	FA1_l6_c31_Cout );

	FA2_l6_c31  : FA 
	PORT MAP ( A =>	PP3(25), B =>	PP4(23), CIN 	=>	PP5(21), S =>	FA2_l6_c31_S, COUT 	=>	FA2_l6_c31_Cout );

	FA3_l6_c31  : FA 
	PORT MAP ( A =>	PP6(19), B =>	PP7(17), CIN 	=>	PP8(15), S =>	FA3_l6_c31_S, COUT 	=>	FA3_l6_c31_Cout );

	HA1_l6_c31  : HA 
	PORT MAP ( A =>	PP9(13), B =>	PP10(11), S =>	HA1_l6_c31_S, COUT 	=>	HA1_l6_c31_Cout );

	FA1_l6_c32  : FA 
	PORT MAP ( A =>	PP0(32), B =>	PP1(30), CIN 	=>	PP2(28), S =>	FA1_l6_c32_S, COUT 	=>	FA1_l6_c32_Cout );

	FA2_l6_c32  : FA 
	PORT MAP ( A =>	PP3(26), B =>	PP4(24), CIN 	=>	PP5(22), S =>	FA2_l6_c32_S, COUT 	=>	FA2_l6_c32_Cout );

	FA3_l6_c32  : FA 
	PORT MAP ( A =>	PP6(20), B =>	PP7(18), CIN 	=>	PP8(16), S =>	FA3_l6_c32_S, COUT 	=>	FA3_l6_c32_Cout );

	FA4_l6_c32  : FA 
	PORT MAP ( A =>	PP9(14), B =>	PP10(12), CIN 	=>	PP11(10), S =>	FA4_l6_c32_S, COUT 	=>	FA4_l6_c32_Cout );

	FA1_l6_c33  : FA 
	PORT MAP ( A =>	PP0(32), B =>	PP1(31), CIN 	=>	PP2(29), S =>	FA1_l6_c33_S, COUT 	=>	FA1_l6_c33_Cout );

	FA2_l6_c33  : FA 
	PORT MAP ( A =>	PP3(27), B =>	PP4(25), CIN 	=>	PP5(23), S =>	FA2_l6_c33_S, COUT 	=>	FA2_l6_c33_Cout );

	FA3_l6_c33  : FA 
	PORT MAP ( A =>	PP6(21), B =>	PP7(19), CIN 	=>	PP8(17), S =>	FA3_l6_c33_S, COUT 	=>	FA3_l6_c33_Cout );

	FA4_l6_c33  : FA 
	PORT MAP ( A =>	PP9(15), B =>	PP10(13), CIN 	=>	PP11(11), S =>	FA4_l6_c33_S, COUT 	=>	FA4_l6_c33_Cout );

	FA1_l6_c34  : FA 
	PORT MAP ( A =>	PP0(32), B =>	PP1(32), CIN 	=>	PP2(30), S =>	FA1_l6_c34_S, COUT 	=>	FA1_l6_c34_Cout );

	FA2_l6_c34  : FA 
	PORT MAP ( A =>	PP3(28), B =>	PP4(26), CIN 	=>	PP5(24), S =>	FA2_l6_c34_S, COUT 	=>	FA2_l6_c34_Cout );

	FA3_l6_c34  : FA 
	PORT MAP ( A =>	PP6(22), B =>	PP7(20), CIN 	=>	PP8(18), S =>	FA3_l6_c34_S, COUT 	=>	FA3_l6_c34_Cout );

	FA4_l6_c34  : FA 
	PORT MAP ( A =>	PP9(16), B =>	PP10(14), CIN 	=>	PP11(12), S =>	FA4_l6_c34_S, COUT 	=>	FA4_l6_c34_Cout );

	FA1_l6_c35  : FA 
	PORT MAP ( A =>	PP0_neg, B =>	PP1_neg, CIN 	=>	PP2(31), S =>	FA1_l6_c35_S, COUT 	=>	FA1_l6_c35_Cout );

	FA2_l6_c35  : FA 
	PORT MAP ( A =>	PP3(29), B =>	PP4(27), CIN 	=>	PP5(25), S =>	FA2_l6_c35_S, COUT 	=>	FA2_l6_c35_Cout );

	FA3_l6_c35  : FA 
	PORT MAP ( A =>	PP6(23), B =>	PP7(21), CIN 	=>	PP8(19), S =>	FA3_l6_c35_S, COUT 	=>	FA3_l6_c35_Cout );

	FA4_l6_c35  : FA 
	PORT MAP ( A =>	PP9(17), B =>	PP10(15), CIN 	=>	PP11(13), S =>	FA4_l6_c35_S, COUT 	=>	FA4_l6_c35_Cout );

	FA1_l6_c36  : FA 
	PORT MAP ( A =>	'1', B =>	PP2(32), CIN 	=>	PP3(30), S =>	FA1_l6_c36_S, COUT 	=>	FA1_l6_c36_Cout );

	FA2_l6_c36  : FA 
	PORT MAP ( A =>	PP4(28), B =>	PP5(26), CIN 	=>	PP6(24), S =>	FA2_l6_c36_S, COUT 	=>	FA2_l6_c36_Cout );

	FA3_l6_c36  : FA 
	PORT MAP ( A =>	PP7(22), B =>	PP8(20), CIN 	=>	PP9(18), S =>	FA3_l6_c36_S, COUT 	=>	FA3_l6_c36_Cout );

	HA1_l6_c36  : HA 
	PORT MAP ( A =>	PP10(16), B =>	PP11(14), S =>	HA1_l6_c36_S, COUT 	=>	HA1_l6_c36_Cout );

	FA1_l6_c37  : FA 
	PORT MAP ( A =>	PP2_neg, B =>	PP3(31), CIN 	=>	PP4(29), S =>	FA1_l6_c37_S, COUT 	=>	FA1_l6_c37_Cout );

	FA2_l6_c37  : FA 
	PORT MAP ( A =>	PP5(27), B =>	PP6(25), CIN 	=>	PP7(23), S =>	FA2_l6_c37_S, COUT 	=>	FA2_l6_c37_Cout );

	FA3_l6_c37  : FA 
	PORT MAP ( A =>	PP8(21), B =>	PP9(19), CIN 	=>	PP10(17), S =>	FA3_l6_c37_S, COUT 	=>	FA3_l6_c37_Cout );

	FA1_l6_c38  : FA 
	PORT MAP ( A =>	'1', B =>	PP3(32), CIN 	=>	PP4(30), S =>	FA1_l6_c38_S, COUT 	=>	FA1_l6_c38_Cout );

	FA2_l6_c38  : FA 
	PORT MAP ( A =>	PP5(28), B =>	PP6(26), CIN 	=>	PP7(24), S =>	FA2_l6_c38_S, COUT 	=>	FA2_l6_c38_Cout );

	HA1_l6_c38  : HA 
	PORT MAP ( A =>	PP8(22), B =>	PP9(20), S =>	HA1_l6_c38_S, COUT 	=>	HA1_l6_c38_Cout );

	FA1_l6_c39  : FA 
	PORT MAP ( A =>	PP3_neg, B =>	PP4(31), CIN 	=>	PP5(29), S =>	FA1_l6_c39_S, COUT 	=>	FA1_l6_c39_Cout );

	FA2_l6_c39  : FA 
	PORT MAP ( A =>	PP6(27), B =>	PP7(25), CIN 	=>	PP8(23), S =>	FA2_l6_c39_S, COUT 	=>	FA2_l6_c39_Cout );

	FA1_l6_c40  : FA 
	PORT MAP ( A =>	'1', B =>	PP4(32), CIN 	=>	PP5(30), S =>	FA1_l6_c40_S, COUT 	=>	FA1_l6_c40_Cout );

	HA1_l6_c40  : HA 
	PORT MAP ( A =>	PP6(28), B =>	PP7(26), S =>	HA1_l6_c40_S, COUT 	=>	HA1_l6_c40_Cout );

	FA1_l6_c41  : FA 
	PORT MAP ( A =>	PP4_neg, B =>	PP5(31), CIN 	=>	PP6(29), S =>	FA1_l6_c41_S, COUT 	=>	FA1_l6_c41_Cout );

	HA1_l6_c42  : HA 
	PORT MAP ( A =>	'1', B =>	PP5(32), S =>	HA1_l6_c42_S, COUT 	=>	HA1_l6_c42_Cout );

	HA1_l5_c16  : HA 
	PORT MAP ( A =>	PP0(16), B =>	PP1(14), S =>	HA1_l5_c16_S, COUT 	=>	HA1_l5_c16_Cout );

	HA1_l5_c17  : HA 
	PORT MAP ( A =>	PP0(17), B =>	PP1(15), S =>	HA1_l5_c17_S, COUT 	=>	HA1_l5_c17_Cout );

	FA1_l5_c18  : FA 
	PORT MAP ( A =>	PP0(18), B =>	PP1(16), CIN 	=>	PP2(14), S =>	FA1_l5_c18_S, COUT 	=>	FA1_l5_c18_Cout );

	HA1_l5_c18  : HA 
	PORT MAP ( A =>	PP3(12), B =>	PP4(10), S =>	HA1_l5_c18_S, COUT 	=>	HA1_l5_c18_Cout );

	FA1_l5_c19  : FA 
	PORT MAP ( A =>	PP0(19), B =>	PP1(17), CIN 	=>	PP2(15), S =>	FA1_l5_c19_S, COUT 	=>	FA1_l5_c19_Cout );

	HA1_l5_c19  : HA 
	PORT MAP ( A =>	PP3(13), B =>	PP4(11), S =>	HA1_l5_c19_S, COUT 	=>	HA1_l5_c19_Cout );

	FA1_l5_c20  : FA 
	PORT MAP ( A =>	PP0(20), B =>	PP1(18), CIN 	=>	PP2(16), S =>	FA1_l5_c20_S, COUT 	=>	FA1_l5_c20_Cout );

	FA2_l5_c20  : FA 
	PORT MAP ( A =>	PP3(14), B =>	PP4(12), CIN 	=>	PP5(10), S =>	FA2_l5_c20_S, COUT 	=>	FA2_l5_c20_Cout );

	HA1_l5_c20  : HA 
	PORT MAP ( A =>	PP6(8), B =>	PP7(6), S =>	HA1_l5_c20_S, COUT 	=>	HA1_l5_c20_Cout );

	FA1_l5_c21  : FA 
	PORT MAP ( A =>	PP0(21), B =>	PP1(19), CIN 	=>	PP2(17), S =>	FA1_l5_c21_S, COUT 	=>	FA1_l5_c21_Cout );

	FA2_l5_c21  : FA 
	PORT MAP ( A =>	PP3(15), B =>	PP4(13), CIN 	=>	PP5(11), S =>	FA2_l5_c21_S, COUT 	=>	FA2_l5_c21_Cout );

	HA1_l5_c21  : HA 
	PORT MAP ( A =>	PP6(9), B =>	PP7(7), S =>	HA1_l5_c21_S, COUT 	=>	HA1_l5_c21_Cout );

	FA1_l5_c22  : FA 
	PORT MAP ( A =>	PP0(22), B =>	PP1(20), CIN 	=>	PP2(18), S =>	FA1_l5_c22_S, COUT 	=>	FA1_l5_c22_Cout );

	FA2_l5_c22  : FA 
	PORT MAP ( A =>	PP3(16), B =>	PP4(14), CIN 	=>	PP5(12), S =>	FA2_l5_c22_S, COUT 	=>	FA2_l5_c22_Cout );

	FA3_l5_c22  : FA 
	PORT MAP ( A =>	PP6(10), B =>	PP7(8), CIN 	=>	PP8(6), S =>	FA3_l5_c22_S, COUT 	=>	FA3_l5_c22_Cout );

	HA1_l5_c22  : HA 
	PORT MAP ( A =>	PP9(4), B =>	PP10(2), S =>	HA1_l5_c22_S, COUT 	=>	HA1_l5_c22_Cout );

	FA1_l5_c23  : FA 
	PORT MAP ( A =>	PP0(23), B =>	PP1(21), CIN 	=>	PP2(19), S =>	FA1_l5_c23_S, COUT 	=>	FA1_l5_c23_Cout );

	FA2_l5_c23  : FA 
	PORT MAP ( A =>	PP3(17), B =>	PP4(15), CIN 	=>	PP5(13), S =>	FA2_l5_c23_S, COUT 	=>	FA2_l5_c23_Cout );

	FA3_l5_c23  : FA 
	PORT MAP ( A =>	PP6(11), B =>	PP7(9), CIN 	=>	PP8(7), S =>	FA3_l5_c23_S, COUT 	=>	FA3_l5_c23_Cout );

	HA1_l5_c23  : HA 
	PORT MAP ( A =>	PP9(5), B =>	PP10(3), S =>	HA1_l5_c23_S, COUT 	=>	HA1_l5_c23_Cout );

	FA1_l5_c24  : FA 
	PORT MAP ( A =>	HA1_l6_c24_S, B =>	PP2(20), CIN 	=>	PP3(18), S =>	FA1_l5_c24_S, COUT 	=>	FA1_l5_c24_Cout );

	FA2_l5_c24  : FA 
	PORT MAP ( A =>	PP4(16), B =>	PP5(14), CIN 	=>	PP6(12), S =>	FA2_l5_c24_S, COUT 	=>	FA2_l5_c24_Cout );

	FA3_l5_c24  : FA 
	PORT MAP ( A =>	PP7(10), B =>	PP8(8), CIN 	=>	PP9(6), S =>	FA3_l5_c24_S, COUT 	=>	FA3_l5_c24_Cout );

	FA4_l5_c24  : FA 
	PORT MAP ( A =>	PP10(4), B =>	PP11(2), CIN 	=>	PP12(0), S =>	FA4_l5_c24_S, COUT 	=>	FA4_l5_c24_Cout );

	FA1_l5_c25  : FA 
	PORT MAP ( A =>	HA1_l6_c24_Cout, B =>	HA1_l6_c25_S, CIN 	=>	PP2(21), S =>	FA1_l5_c25_S, COUT 	=>	FA1_l5_c25_Cout );

	FA2_l5_c25  : FA 
	PORT MAP ( A =>	PP3(19), B =>	PP4(17), CIN 	=>	PP5(15), S =>	FA2_l5_c25_S, COUT 	=>	FA2_l5_c25_Cout );

	FA3_l5_c25  : FA 
	PORT MAP ( A =>	PP6(13), B =>	PP7(11), CIN 	=>	PP8(9), S =>	FA3_l5_c25_S, COUT 	=>	FA3_l5_c25_Cout );

	FA4_l5_c25  : FA 
	PORT MAP ( A =>	PP9(7), B =>	PP10(5), CIN 	=>	PP11(3), S =>	FA4_l5_c25_S, COUT 	=>	FA4_l5_c25_Cout );

	FA1_l5_c26  : FA 
	PORT MAP ( A =>	HA1_l6_c25_Cout, B =>	HA1_l6_c26_S, CIN 	=>	FA1_l6_c26_S, S =>	FA1_l5_c26_S, COUT 	=>	FA1_l5_c26_Cout );

	FA2_l5_c26  : FA 
	PORT MAP ( A =>	PP5(16), B =>	PP6(14), CIN 	=>	PP7(12), S =>	FA2_l5_c26_S, COUT 	=>	FA2_l5_c26_Cout );

	FA3_l5_c26  : FA 
	PORT MAP ( A =>	PP8(10), B =>	PP9(8), CIN 	=>	PP10(6), S =>	FA3_l5_c26_S, COUT 	=>	FA3_l5_c26_Cout );

	FA4_l5_c26  : FA 
	PORT MAP ( A =>	PP11(4), B =>	PP12(2), CIN 	=>	PP13(0), S =>	FA4_l5_c26_S, COUT 	=>	FA4_l5_c26_Cout );

	FA1_l5_c27  : FA 
	PORT MAP ( A =>	HA1_l6_c26_Cout, B =>	FA1_l6_c26_Cout, CIN 	=>	HA1_l6_c27_S, S =>	FA1_l5_c27_S, COUT 	=>	FA1_l5_c27_Cout );

	FA2_l5_c27  : FA 
	PORT MAP ( A =>	FA1_l6_c27_S, B =>	PP5(17), CIN 	=>	PP6(15), S =>	FA2_l5_c27_S, COUT 	=>	FA2_l5_c27_Cout );

	FA3_l5_c27  : FA 
	PORT MAP ( A =>	PP7(13), B =>	PP8(11), CIN 	=>	PP9(9), S =>	FA3_l5_c27_S, COUT 	=>	FA3_l5_c27_Cout );

	FA4_l5_c27  : FA 
	PORT MAP ( A =>	PP10(7), B =>	PP11(5), CIN 	=>	PP12(3), S =>	FA4_l5_c27_S, COUT 	=>	FA4_l5_c27_Cout );

	FA1_l5_c28  : FA 
	PORT MAP ( A =>	HA1_l6_c27_Cout, B =>	FA1_l6_c27_Cout, CIN 	=>	HA1_l6_c28_S, S =>	FA1_l5_c28_S, COUT 	=>	FA1_l5_c28_Cout );

	FA2_l5_c28  : FA 
	PORT MAP ( A =>	FA2_l6_c28_S, B =>	FA1_l6_c28_S, CIN 	=>	PP8(12), S =>	FA2_l5_c28_S, COUT 	=>	FA2_l5_c28_Cout );

	FA3_l5_c28  : FA 
	PORT MAP ( A =>	PP9(10), B =>	PP10(8), CIN 	=>	PP11(6), S =>	FA3_l5_c28_S, COUT 	=>	FA3_l5_c28_Cout );

	FA4_l5_c28  : FA 
	PORT MAP ( A =>	PP12(4), B =>	PP13(2), CIN 	=>	PP14(0), S =>	FA4_l5_c28_S, COUT 	=>	FA4_l5_c28_Cout );

	
	FA1_l5_c29  : FA 
	PORT MAP ( A =>	HA1_l6_c28_Cout, B =>	FA2_l6_c28_Cout, CIN 	=>	FA1_l6_c28_Cout, S =>	FA1_l5_c29_S, COUT 	=>	FA1_l5_c29_Cout );

	FA2_l5_c29  : FA 
	PORT MAP ( A =>	HA1_l6_c29_S, B =>	FA2_l6_c29_S, CIN 	=>	FA1_l6_c29_S, S =>	FA2_l5_c29_S, COUT 	=>	FA2_l5_c29_Cout );

	FA3_l5_c29  : FA 
	PORT MAP ( A =>	PP8(13), B =>	PP9(11), CIN 	=>	PP10(9), S =>	FA3_l5_c29_S, COUT 	=>	FA3_l5_c29_Cout );

	FA4_l5_c29  : FA 
	PORT MAP ( A =>	PP11(7), B =>	PP12(5), CIN 	=>	PP13(3), S =>	FA4_l5_c29_S, COUT 	=>	FA4_l5_c29_Cout );

	FA1_l5_c30  : FA 
	PORT MAP ( A =>	HA1_l6_c29_Cout, B =>	FA2_l6_c29_Cout, CIN 	=>	FA1_l6_c29_Cout, S =>	FA1_l5_c30_S, COUT 	=>	FA1_l5_c30_Cout );

	FA2_l5_c30  : FA 
	PORT MAP ( A =>	HA1_l6_c30_S, B =>	FA3_l6_c30_S, CIN 	=>	FA2_l6_c30_S, S =>	FA2_l5_c30_S, COUT 	=>	FA2_l5_c30_Cout );

	FA3_l5_c30  : FA 
	PORT MAP ( A =>	FA1_l6_c30_S, B =>	PP11(8), CIN 	=>	PP12(6), S =>	FA3_l5_c30_S, COUT 	=>	FA3_l5_c30_Cout );

	FA4_l5_c30  : FA 
	PORT MAP ( A =>	PP13(4), B =>	PP14(2), CIN 	=>	PP15(0), S =>	FA4_l5_c30_S, COUT 	=>	FA4_l5_c30_Cout );

	FA1_l5_c31  : FA 
	PORT MAP ( A =>	HA1_l6_c30_Cout, B =>	FA3_l6_c30_Cout, CIN 	=>	FA2_l6_c30_Cout, S =>	FA1_l5_c31_S, COUT 	=>	FA1_l5_c31_Cout );

	FA2_l5_c31  : FA 
	PORT MAP ( A =>	FA1_l6_c30_Cout, B =>	HA1_l6_c31_S, CIN 	=>	FA3_l6_c31_S, S =>	FA2_l5_c31_S, COUT 	=>	FA2_l5_c31_Cout );

	FA3_l5_c31  : FA 
	PORT MAP ( A =>	FA2_l6_c31_S, B =>	FA1_l6_c31_S, CIN 	=>	PP11(9), S =>	FA3_l5_c31_S, COUT 	=>	FA3_l5_c31_Cout );

	FA4_l5_c31  : FA 
	PORT MAP ( A =>	PP12(7), B =>	PP13(5), CIN 	=>	PP14(3), S =>	FA4_l5_c31_S, COUT 	=>	FA4_l5_c31_Cout );

	FA1_l5_c32  : FA 
	PORT MAP ( A =>	HA1_l6_c31_Cout, B =>	FA3_l6_c31_Cout, CIN 	=>	FA2_l6_c31_Cout, S =>	FA1_l5_c32_S, COUT 	=>	FA1_l5_c32_Cout );

	FA2_l5_c32  : FA 
	PORT MAP ( A =>	FA1_l6_c31_Cout, B =>	FA4_l6_c32_S, CIN 	=>	FA3_l6_c32_S, S =>	FA2_l5_c32_S, COUT 	=>	FA2_l5_c32_Cout );

	FA3_l5_c32  : FA 
	PORT MAP ( A =>	FA2_l6_c32_S, B =>	FA1_l6_c32_S, CIN 	=>	PP12(8), S =>	FA3_l5_c32_S, COUT 	=>	FA3_l5_c32_Cout );

	FA4_l5_c32  : FA 
	PORT MAP ( A =>	PP13(6), B =>	PP14(4), CIN 	=>	PP15(2), S =>	FA4_l5_c32_S, COUT 	=>	FA4_l5_c32_Cout );

	FA1_l5_c33  : FA 
	PORT MAP ( A =>	FA4_l6_c32_Cout, B =>	FA3_l6_c32_Cout, CIN 	=>	FA2_l6_c32_Cout, S =>	FA1_l5_c33_S, COUT 	=>	FA1_l5_c33_Cout );

	FA2_l5_c33  : FA 
	PORT MAP ( A =>	FA1_l6_c32_Cout, B =>	FA4_l6_c33_S, CIN 	=>	FA3_l6_c33_S, S =>	FA2_l5_c33_S, COUT 	=>	FA2_l5_c33_Cout );

	FA3_l5_c33  : FA 
	PORT MAP ( A =>	FA2_l6_c33_S, B =>	FA1_l6_c33_S, CIN 	=>	PP12(9), S =>	FA3_l5_c33_S, COUT 	=>	FA3_l5_c33_Cout );

	FA4_l5_c33  : FA 
	PORT MAP ( A =>	PP13(7), B =>	PP14(5), CIN 	=>	PP15(3), S =>	FA4_l5_c33_S, COUT 	=>	FA4_l5_c33_Cout );

	FA1_l5_c34  : FA 
	PORT MAP ( A =>	FA4_l6_c33_Cout, B =>	FA3_l6_c33_Cout, CIN 	=>	FA2_l6_c33_Cout, S =>	FA1_l5_c34_S, COUT 	=>	FA1_l5_c34_Cout );

	FA2_l5_c34  : FA 
	PORT MAP ( A =>	FA1_l6_c33_Cout, B =>	FA4_l6_c34_S, CIN 	=>	FA3_l6_c34_S, S =>	FA2_l5_c34_S, COUT 	=>	FA2_l5_c34_Cout );

	FA3_l5_c34  : FA 
	PORT MAP ( A =>	FA2_l6_c34_S, B =>	FA1_l6_c34_S, CIN 	=>	PP12(10), S =>	FA3_l5_c34_S, COUT 	=>	FA3_l5_c34_Cout );

	FA4_l5_c34  : FA 
	PORT MAP ( A =>	PP13(8), B =>	PP14(6), CIN 	=>	PP15(4), S =>	FA4_l5_c34_S, COUT 	=>	FA4_l5_c34_Cout );

	FA1_l5_c35  : FA 
	PORT MAP ( A =>	FA4_l6_c34_Cout, B =>	FA3_l6_c34_Cout, CIN 	=>	FA2_l6_c34_Cout, S =>	FA1_l5_c35_S, COUT 	=>	FA1_l5_c35_Cout );

	FA2_l5_c35  : FA 
	PORT MAP ( A =>	FA1_l6_c34_Cout, B =>	FA4_l6_c35_S, CIN 	=>	FA3_l6_c35_S, S =>	FA2_l5_c35_S, COUT 	=>	FA2_l5_c35_Cout );

	FA3_l5_c35  : FA 
	PORT MAP ( A =>	FA2_l6_c35_S, B =>	FA1_l6_c35_S, CIN 	=>	PP12(11), S =>	FA3_l5_c35_S, COUT 	=>	FA3_l5_c35_Cout );

	FA4_l5_c35  : FA 
	PORT MAP ( A =>	PP13(9), B =>	PP14(7), CIN 	=>	PP15(5), S =>	FA4_l5_c35_S, COUT 	=>	FA4_l5_c35_Cout );

	FA1_l5_c36  : FA 
	PORT MAP ( A =>	FA4_l6_c35_Cout, B =>	FA3_l6_c35_Cout, CIN 	=>	FA2_l6_c35_Cout, S =>	FA1_l5_c36_S, COUT 	=>	FA1_l5_c36_Cout );

	FA2_l5_c36  : FA 
	PORT MAP ( A =>	FA1_l6_c35_Cout, B =>	HA1_l6_c36_S, CIN 	=>	FA3_l6_c36_S, S =>	FA2_l5_c36_S, COUT 	=>	FA2_l5_c36_Cout );

	FA3_l5_c36  : FA 
	PORT MAP ( A =>	FA2_l6_c36_S, B =>	FA1_l6_c36_S, CIN 	=>	PP12(12), S =>	FA3_l5_c36_S, COUT 	=>	FA3_l5_c36_Cout );

	FA4_l5_c36  : FA 
	PORT MAP ( A =>	PP13(10), B =>	PP14(8), CIN 	=>	PP15(6), S =>	FA4_l5_c36_S, COUT 	=>	FA4_l5_c36_Cout );

	FA1_l5_c37  : FA 
	PORT MAP ( A =>	HA1_l6_c36_Cout, B =>	FA3_l6_c36_Cout, CIN 	=>	FA2_l6_c36_Cout, S =>	FA1_l5_c37_S, COUT 	=>	FA1_l5_c37_Cout );

	FA2_l5_c37  : FA 
	PORT MAP ( A =>	FA1_l6_c36_Cout, B =>	FA3_l6_c37_S, CIN 	=>	FA2_l6_c37_S, S =>	FA2_l5_c37_S, COUT 	=>	FA2_l5_c37_Cout );

	FA3_l5_c37  : FA 
	PORT MAP ( A =>	FA1_l6_c37_S, B =>	PP11(15), CIN 	=>	PP12(13), S =>	FA3_l5_c37_S, COUT 	=>	FA3_l5_c37_Cout );

	FA4_l5_c37  : FA 
	PORT MAP ( A =>	PP13(11), B =>	PP14(9), CIN 	=>	PP15(7), S =>	FA4_l5_c37_S, COUT 	=>	FA4_l5_c37_Cout );

	FA1_l5_c38  : FA 
	PORT MAP ( A =>	FA3_l6_c37_Cout, B =>	FA2_l6_c37_Cout, CIN 	=>	FA1_l6_c37_Cout, S =>	FA1_l5_c38_S, COUT 	=>	FA1_l5_c38_Cout );

	FA2_l5_c38  : FA 
	PORT MAP ( A =>	HA1_l6_c38_S, B =>	FA2_l6_c38_S, CIN 	=>	FA1_l6_c38_S, S =>	FA2_l5_c38_S, COUT 	=>	FA2_l5_c38_Cout );

	FA3_l5_c38  : FA 
	PORT MAP ( A =>	PP10(18), B =>	PP11(16), CIN 	=>	PP12(14), S =>	FA3_l5_c38_S, COUT 	=>	FA3_l5_c38_Cout );

	FA4_l5_c38  : FA 
	PORT MAP ( A =>	PP13(12), B =>	PP14(10), CIN 	=>	PP15(8), S =>	FA4_l5_c38_S, COUT 	=>	FA4_l5_c38_Cout );

	FA1_l5_c39  : FA 
	PORT MAP ( A =>	HA1_l6_c38_Cout, B =>	FA2_l6_c38_Cout, CIN 	=>	FA1_l6_c38_Cout, S =>	FA1_l5_c39_S, COUT 	=>	FA1_l5_c39_Cout );

	FA2_l5_c39  : FA 
	PORT MAP ( A =>	FA2_l6_c39_S, B =>	FA1_l6_c39_S, CIN 	=>	PP9(21), S =>	FA2_l5_c39_S, COUT 	=>	FA2_l5_c39_Cout );

	FA3_l5_c39  : FA 
	PORT MAP ( A =>	PP10(19), B =>	PP11(17), CIN 	=>	PP12(15), S =>	FA3_l5_c39_S, COUT 	=>	FA3_l5_c39_Cout );

	FA4_l5_c39  : FA 
	PORT MAP ( A =>	PP13(13), B =>	PP14(11), CIN 	=>	PP15(9), S =>	FA4_l5_c39_S, COUT 	=>	FA4_l5_c39_Cout );

	FA1_l5_c40  : FA 
	PORT MAP ( A =>	FA2_l6_c39_Cout, B =>	FA1_l6_c39_Cout, CIN 	=>	HA1_l6_c40_S, S =>	FA1_l5_c40_S, COUT 	=>	FA1_l5_c40_Cout );

	FA2_l5_c40  : FA 
	PORT MAP ( A =>	FA1_l6_c40_S, B =>	PP8(24), CIN 	=>	PP9(22), S =>	FA2_l5_c40_S, COUT 	=>	FA2_l5_c40_Cout );

	FA3_l5_c40  : FA 
	PORT MAP ( A =>	PP10(20), B =>	PP11(18), CIN 	=>	PP12(16), S =>	FA3_l5_c40_S, COUT 	=>	FA3_l5_c40_Cout );

	FA4_l5_c40  : FA 
	PORT MAP ( A =>	PP13(14), B =>	PP14(12), CIN 	=>	PP15(10), S =>	FA4_l5_c40_S, COUT 	=>	FA4_l5_c40_Cout );

	FA1_l5_c41  : FA 
	PORT MAP ( A =>	HA1_l6_c40_Cout, B =>	FA1_l6_c40_Cout, CIN 	=>	FA1_l6_c41_S, S =>	FA1_l5_c41_S, COUT 	=>	FA1_l5_c41_Cout );

	FA2_l5_c41  : FA 
	PORT MAP ( A =>	PP7(27), B =>	PP8(25), CIN 	=>	PP9(23), S =>	FA2_l5_c41_S, COUT 	=>	FA2_l5_c41_Cout );

	FA3_l5_c41  : FA 
	PORT MAP ( A =>	PP10(21), B =>	PP11(19), CIN 	=>	PP12(17), S =>	FA3_l5_c41_S, COUT 	=>	FA3_l5_c41_Cout );

	FA4_l5_c41  : FA 
	PORT MAP ( A =>	PP13(15), B =>	PP14(13), CIN 	=>	PP15(11), S =>	FA4_l5_c41_S, COUT 	=>	FA4_l5_c41_Cout );

	FA1_l5_c42  : FA 
	PORT MAP ( A =>	FA1_l6_c41_Cout, B =>	HA1_l6_c42_S, CIN 	=>	PP6(30), S =>	FA1_l5_c42_S, COUT 	=>	FA1_l5_c42_Cout );

	FA2_l5_c42  : FA 
	PORT MAP ( A =>	PP7(28), B =>	PP8(26), CIN 	=>	PP9(24), S =>	FA2_l5_c42_S, COUT 	=>	FA2_l5_c42_Cout );

	FA3_l5_c42  : FA 
	PORT MAP ( A =>	PP10(22), B =>	PP11(20), CIN 	=>	PP12(18), S =>	FA3_l5_c42_S, COUT 	=>	FA3_l5_c42_Cout );

	FA4_l5_c42  : FA 
	PORT MAP ( A =>	PP13(16), B =>	PP14(14), CIN 	=>	PP15(12), S =>	FA4_l5_c42_S, COUT 	=>	FA4_l5_c42_Cout );

	FA1_l5_c43  : FA 
	PORT MAP ( A =>	HA1_l6_c42_Cout, B =>	PP5_neg, CIN 	=>	PP6(31), S =>	FA1_l5_c43_S, COUT 	=>	FA1_l5_c43_Cout );

	FA2_l5_c43  : FA 
	PORT MAP ( A =>	PP7(29), B =>	PP8(27), CIN 	=>	PP9(25), S =>	FA2_l5_c43_S, COUT 	=>	FA2_l5_c43_Cout );

	FA3_l5_c43  : FA 
	PORT MAP ( A =>	PP10(23), B =>	PP11(21), CIN 	=>	PP12(19), S =>	FA3_l5_c43_S, COUT 	=>	FA3_l5_c43_Cout );

	FA4_l5_c43  : FA 
	PORT MAP ( A =>	PP13(17), B =>	PP14(15), CIN 	=>	PP15(13), S =>	FA4_l5_c43_S, COUT 	=>	FA4_l5_c43_Cout );

	FA1_l5_c44  : FA 
	PORT MAP ( A =>	'1', B =>	PP6(32), CIN 	=>	PP7(30), S =>	FA1_l5_c44_S, COUT 	=>	FA1_l5_c44_Cout );

	FA2_l5_c44  : FA 
	PORT MAP ( A =>	PP8(28), B =>	PP9(26), CIN 	=>	PP10(24), S =>	FA2_l5_c44_S, COUT 	=>	FA2_l5_c44_Cout );

	FA3_l5_c44  : FA 
	PORT MAP ( A =>	PP11(22), B =>	PP12(20), CIN 	=>	PP13(18), S =>	FA3_l5_c44_S, COUT 	=>	FA3_l5_c44_Cout );

	HA1_l5_c44  : HA 
	PORT MAP ( A =>	PP14(16), B =>	PP15(14), S =>	HA1_l5_c44_S, COUT 	=>	HA1_l5_c44_Cout );

	FA1_l5_c45  : FA 
	PORT MAP ( A =>	PP6_neg, B =>	PP7(31), CIN 	=>	PP8(29), S =>	FA1_l5_c45_S, COUT 	=>	FA1_l5_c45_Cout );

	FA2_l5_c45  : FA 
	PORT MAP ( A =>	PP9(27), B =>	PP10(25), CIN 	=>	PP11(23), S =>	FA2_l5_c45_S, COUT 	=>	FA2_l5_c45_Cout );

	FA3_l5_c45  : FA
	PORT MAP ( A =>	PP12(21), B =>	PP13(19), CIN 	=>	PP14(17), S =>	FA3_l5_c45_S, COUT 	=>	FA3_l5_c45_Cout );

	FA1_l5_c46  : FA 
	PORT MAP ( A =>	'1', B =>	PP7(32), CIN 	=>	PP8(30), S =>	FA1_l5_c46_S, COUT 	=>	FA1_l5_c46_Cout );

	FA2_l5_c46  : FA 
	PORT MAP ( A =>	PP9(28), B =>	PP10(26), CIN 	=>	PP11(24), S =>	FA2_l5_c46_S, COUT 	=>	FA2_l5_c46_Cout );

	HA1_l5_c46  : HA 
	PORT MAP ( A =>	PP12(22), B =>	PP13(20), S =>	HA1_l5_c46_S, COUT 	=>	HA1_l5_c46_Cout );

	FA1_l5_c47  : FA 
	PORT MAP ( A =>	PP7_neg, B =>	PP8(31), CIN 	=>	PP9(29), S =>	FA1_l5_c47_S, COUT 	=>	FA1_l5_c47_Cout );

	FA2_l5_c47  : FA 
	PORT MAP ( A =>	PP10(27), B =>	PP11(25), CIN 	=>	PP12(23), S =>	FA2_l5_c47_S, COUT 	=>	FA2_l5_c47_Cout );

	FA1_l5_c48  : FA 
	PORT MAP ( A =>	'1', B =>	PP8(32), CIN 	=>	PP9(30), S =>	FA1_l5_c48_S, COUT 	=>	FA1_l5_c48_Cout );

	HA1_l5_c48  : HA 
	PORT MAP ( A =>	PP10(28), B =>	PP11(26), S =>	HA1_l5_c48_S, COUT 	=>	HA1_l5_c48_Cout );

	FA1_l5_c49  : FA 
	PORT MAP ( A =>	PP8_neg, B =>	PP9(31), CIN 	=>	PP10(29), S =>	FA1_l5_c49_S, COUT 	=>	FA1_l5_c49_Cout );

	HA1_l5_c50  : HA 
	PORT MAP ( A =>	'1', B =>	PP9(32), S =>	HA1_l5_c50_S, COUT 	=>	HA1_l5_c50_Cout );

	HA1_l4_c10  : HA 
	PORT MAP ( A =>	PP0(10), B =>	PP1(8), S =>	HA1_l4_c10_S, COUT 	=>	HA1_l4_c10_Cout );

	HA1_l4_c11  : HA 
	PORT MAP ( A =>	PP0(11), B =>	PP1(9), S =>	HA1_l4_c11_S, COUT 	=>	HA1_l4_c11_Cout );

	FA1_l4_c12  : FA 
	PORT MAP ( A =>	PP0(12), B =>	PP1(10), CIN 	=>	PP2(8), S =>	FA1_l4_c12_S, COUT 	=>	FA1_l4_c12_Cout );

	HA1_l4_c12  : HA 
	PORT MAP ( A =>	PP3(6), B =>	PP4(4), S =>	HA1_l4_c12_S, COUT 	=>	HA1_l4_c12_Cout );

	FA1_l4_c13  : FA 
	PORT MAP ( A =>	PP0(13), B =>	PP1(11), CIN 	=>	PP2(9), S =>	FA1_l4_c13_S, COUT 	=>	FA1_l4_c13_Cout );

	HA1_l4_c13  : HA 
	PORT MAP ( A =>	PP3(7), B =>	PP4(5), S =>	HA1_l4_c13_S, COUT 	=>	HA1_l4_c13_Cout );

	FA1_l4_c14  : FA 
	PORT MAP ( A =>	PP0(14), B =>	PP1(12), CIN 	=>	PP2(10), S =>	FA1_l4_c14_S, COUT 	=>	FA1_l4_c14_Cout );

	FA2_l4_c14  : FA 
	PORT MAP ( A =>	PP3(8), B =>	PP4(6), CIN 	=>	PP5(4), S =>	FA2_l4_c14_S, COUT 	=>	FA2_l4_c14_Cout );

	HA1_l4_c14  : HA 
	PORT MAP ( A =>	PP6(2), B =>	PP7(0), S =>	HA1_l4_c14_S, COUT 	=>	HA1_l4_c14_Cout );

	FA1_l4_c15  : FA 
	PORT MAP ( A =>	PP0(15), B =>	PP1(13), CIN 	=>	PP2(11), S =>	FA1_l4_c15_S, COUT 	=>	FA1_l4_c15_Cout );

	FA2_l4_c15  : FA 
	PORT MAP ( A =>	PP3(9), B =>	PP4(7), CIN 	=>	PP5(5), S =>	FA2_l4_c15_S, COUT 	=>	FA2_l4_c15_Cout );

	HA1_l4_c15  : HA 
	PORT MAP ( A =>	PP6(3), B =>	PP7(1), S =>	HA1_l4_c15_S, COUT 	=>	HA1_l4_c15_Cout );

	FA1_l4_c16  : FA 
	PORT MAP ( A =>	HA1_l5_c16_S, B =>	PP2(12), CIN 	=>	PP3(10), S =>	FA1_l4_c16_S, COUT 	=>	FA1_l4_c16_Cout );

	FA2_l4_c16  : FA 
	PORT MAP ( A =>	PP4(8), B =>	PP5(6), CIN 	=>	PP6(4), S =>	FA2_l4_c16_S, COUT 	=>	FA2_l4_c16_Cout );

	FA3_l4_c16  : FA 
	PORT MAP ( A =>	PP7(2), B =>	PP8(0), CIN 	=>	PP8(32), S =>	FA3_l4_c16_S, COUT 	=>	FA3_l4_c16_Cout );

	FA1_l4_c17  : FA 
	PORT MAP ( A =>	HA1_l5_c16_Cout, B =>	HA1_l5_c17_S, CIN 	=>	PP2(13), S =>	FA1_l4_c17_S, COUT 	=>	FA1_l4_c17_Cout );

	FA2_l4_c17  : FA 
	PORT MAP ( A =>	PP3(11), B =>	PP4(9), CIN 	=>	PP5(7), S =>	FA2_l4_c17_S, COUT 	=>	FA2_l4_c17_Cout );

	FA3_l4_c17  : FA 
	PORT MAP ( A =>	PP6(5), B =>	PP7(3), CIN 	=>	PP8(1), S =>	FA3_l4_c17_S, COUT 	=>	FA3_l4_c17_Cout );

	FA1_l4_c18  : FA 
	PORT MAP ( A =>	HA1_l5_c17_Cout, B =>	HA1_l5_c18_S, CIN 	=>	FA1_l5_c18_S, S =>	FA1_l4_c18_S, COUT 	=>	FA1_l4_c18_Cout );

	FA2_l4_c18  : FA 
	PORT MAP ( A =>	PP5(8), B =>	PP6(6), CIN 	=>	PP7(4), S =>	FA2_l4_c18_S, COUT 	=>	FA2_l4_c18_Cout );

	FA3_l4_c18  : FA 
	PORT MAP ( A =>	PP8(2), B =>	PP9(0), CIN 	=>	PP9(32), S =>	FA3_l4_c18_S, COUT 	=>	FA3_l4_c18_Cout );

	FA1_l4_c19  : FA 
	PORT MAP ( A =>	HA1_l5_c18_Cout, B =>	FA1_l5_c18_Cout, CIN 	=>	HA1_l5_c19_S, S =>	FA1_l4_c19_S, COUT 	=>	FA1_l4_c19_Cout );

	FA2_l4_c19  : FA 
	PORT MAP ( A =>	FA1_l5_c19_S, B =>	PP5(9), CIN 	=>	PP6(7), S =>	FA2_l4_c19_S, COUT 	=>	FA2_l4_c19_Cout );

	FA3_l4_c19  : FA 
	PORT MAP ( A =>	PP7(5), B =>	PP8(3), CIN 	=>	PP9(1), S =>	FA3_l4_c19_S, COUT 	=>	FA3_l4_c19_Cout );

	FA1_l4_c20  : FA 
	PORT MAP ( A =>	HA1_l5_c19_Cout, B =>	FA1_l5_c19_Cout, CIN 	=>	HA1_l5_c20_S, S =>	FA1_l4_c20_S, COUT 	=>	FA1_l4_c20_Cout );

	FA2_l4_c20  : FA 
	PORT MAP ( A =>	FA2_l5_c20_S, B =>	FA1_l5_c20_S, CIN 	=>	PP8(4), S =>	FA2_l4_c20_S, COUT 	=>	FA2_l4_c20_Cout );

	FA3_l4_c20  : FA 
	PORT MAP ( A =>	PP9(2), B =>	PP10(0), CIN 	=>	PP10(32), S =>	FA3_l4_c20_S, COUT 	=>	FA3_l4_c20_Cout );

	FA1_l4_c21  : FA 
	PORT MAP ( A =>	HA1_l5_c20_Cout, B =>	FA2_l5_c20_Cout, CIN 	=>	FA1_l5_c20_Cout, S =>	FA1_l4_c21_S, COUT 	=>	FA1_l4_c21_Cout );

	FA2_l4_c21  : FA 
	PORT MAP ( A =>	HA1_l5_c21_S, B =>	FA2_l5_c21_S, CIN 	=>	FA1_l5_c21_S, S =>	FA2_l4_c21_S, COUT 	=>	FA2_l4_c21_Cout );

	FA3_l4_c21  : FA 
	PORT MAP ( A =>	PP8(5), B =>	PP9(3), CIN 	=>	PP10(1), S =>	FA3_l4_c21_S, COUT 	=>	FA3_l4_c21_Cout );

	FA1_l4_c22  : FA 
	PORT MAP ( A =>	HA1_l5_c21_Cout, B =>	FA2_l5_c21_Cout, CIN 	=>	FA1_l5_c21_Cout, S =>	FA1_l4_c22_S, COUT 	=>	FA1_l4_c22_Cout );

	FA2_l4_c22  : FA 
	PORT MAP ( A =>	HA1_l5_c22_S, B =>	FA3_l5_c22_S, CIN 	=>	FA2_l5_c22_S, S =>	FA2_l4_c22_S, COUT 	=>	FA2_l4_c22_Cout );

	FA3_l4_c22  : FA 
	PORT MAP ( A =>	FA1_l5_c22_S, B =>	PP11(0), CIN 	=>	PP11(32), S =>	FA3_l4_c22_S, COUT 	=>	FA3_l4_c22_Cout );

	FA1_l4_c23  : FA 
	PORT MAP ( A =>	HA1_l5_c22_Cout, B =>	FA3_l5_c22_Cout, CIN 	=>	FA2_l5_c22_Cout, S =>	FA1_l4_c23_S, COUT 	=>	FA1_l4_c23_Cout );

	FA2_l4_c23  : FA 
	PORT MAP ( A =>	FA1_l5_c22_Cout, B =>	HA1_l5_c23_S, CIN 	=>	FA3_l5_c23_S, S =>	FA2_l4_c23_S, COUT 	=>	FA2_l4_c23_Cout );

	FA3_l4_c23  : FA 
	PORT MAP ( A =>	FA2_l5_c23_S, B =>	FA1_l5_c23_S, CIN 	=>	PP11(1), S =>	FA3_l4_c23_S, COUT 	=>	FA3_l4_c23_Cout );

	FA1_l4_c24  : FA 
	PORT MAP ( A =>	HA1_l5_c23_Cout, B =>	FA3_l5_c23_Cout, CIN 	=>	FA2_l5_c23_Cout, S =>	FA1_l4_c24_S, COUT 	=>	FA1_l4_c24_Cout );

	FA2_l4_c24  : FA 
	PORT MAP ( A =>	FA1_l5_c23_Cout, B =>	FA4_l5_c24_S, CIN 	=>	FA3_l5_c24_S, S =>	FA2_l4_c24_S, COUT 	=>	FA2_l4_c24_Cout );

	FA3_l4_c24  : FA 
	PORT MAP ( A =>	FA2_l5_c24_S, B =>	FA1_l5_c24_S, CIN 	=>	PP12(32), S =>	FA3_l4_c24_S, COUT 	=>	FA3_l4_c24_Cout );

	FA1_l4_c25  : FA 
	PORT MAP ( A =>	FA4_l5_c24_Cout, B =>	FA3_l5_c24_Cout, CIN 	=>	FA2_l5_c24_Cout, S =>	FA1_l4_c25_S, COUT 	=>	FA1_l4_c25_Cout );

	FA2_l4_c25  : FA 
	PORT MAP ( A =>	FA1_l5_c24_Cout, B =>	FA4_l5_c25_S, CIN 	=>	FA3_l5_c25_S, S =>	FA2_l4_c25_S, COUT 	=>	FA2_l4_c25_Cout );

	FA3_l4_c25  : FA 
	PORT MAP ( A =>	FA2_l5_c25_S, B =>	FA1_l5_c25_S, CIN 	=>	PP12(1), S =>	FA3_l4_c25_S, COUT 	=>	FA3_l4_c25_Cout );

	FA1_l4_c26  : FA
	PORT MAP ( A =>	FA4_l5_c25_Cout, B =>	FA3_l5_c25_Cout, CIN 	=>	FA2_l5_c25_Cout, S =>	FA1_l4_c26_S, COUT 	=>	FA1_l4_c26_Cout );

	FA2_l4_c26  : FA
	PORT MAP ( A =>	FA1_l5_c25_Cout, B =>	FA4_l5_c26_S, CIN 	=>	FA3_l5_c26_S, S =>	FA2_l4_c26_S, COUT 	=>	FA2_l4_c26_Cout );

	FA3_l4_c26  : FA
	PORT MAP ( A =>	FA2_l5_c26_S, B =>	FA1_l5_c26_S, CIN 	=>	PP13(32), S =>	FA3_l4_c26_S, COUT 	=>	FA3_l4_c26_Cout );

	FA1_l4_c27  : FA 
	PORT MAP ( A =>	FA4_l5_c26_Cout, B =>	FA3_l5_c26_Cout, CIN 	=>	FA2_l5_c26_Cout, S =>	FA1_l4_c27_S, COUT 	=>	FA1_l4_c27_Cout );

	FA2_l4_c27  : FA
	PORT MAP ( A =>	FA1_l5_c26_Cout, B =>	FA4_l5_c27_S, CIN 	=>	FA3_l5_c27_S, S =>	FA2_l4_c27_S, COUT 	=>	FA2_l4_c27_Cout );

	FA3_l4_c27  : FA 
	PORT MAP ( A =>	FA2_l5_c27_S, B =>	FA1_l5_c27_S, CIN 	=>	PP13(1), S =>	FA3_l4_c27_S, COUT 	=>	FA3_l4_c27_Cout );

	FA1_l4_c28  : FA 
	PORT MAP ( A =>	FA4_l5_c27_Cout, B =>	FA3_l5_c27_Cout, CIN 	=>	FA2_l5_c27_Cout, S =>	FA1_l4_c28_S, COUT 	=>	FA1_l4_c28_Cout );

	FA2_l4_c28  : FA 
	PORT MAP ( A =>	FA1_l5_c27_Cout, B =>	FA4_l5_c28_S, CIN 	=>	FA3_l5_c28_S, S =>	FA2_l4_c28_S, COUT 	=>	FA2_l4_c28_Cout );

	FA3_l4_c28  : FA 
	PORT MAP ( A =>	FA2_l5_c28_S, B =>	FA1_l5_c28_S, CIN 	=>	PP14(32), S =>	FA3_l4_c28_S, COUT 	=>	FA3_l4_c28_Cout );

	FA1_l4_c29  : FA 
	PORT MAP ( A =>	FA4_l5_c28_Cout, B =>	FA3_l5_c28_Cout, CIN 	=>	FA2_l5_c28_Cout, S =>	FA1_l4_c29_S, COUT 	=>	FA1_l4_c29_Cout );

	FA2_l4_c29  : FA 
	PORT MAP ( A =>	FA1_l5_c28_Cout, B =>	FA4_l5_c29_S, CIN 	=>	FA3_l5_c29_S, S =>	FA2_l4_c29_S, COUT 	=>	FA2_l4_c29_Cout );

	FA3_l4_c29  : FA 
	PORT MAP ( A =>	FA2_l5_c29_S, B =>	FA1_l5_c29_S, CIN 	=>	PP14(1), S =>	FA3_l4_c29_S, COUT 	=>	FA3_l4_c29_Cout );

	FA1_l4_c30  : FA 
	PORT MAP ( A =>	FA4_l5_c29_Cout, B =>	FA3_l5_c29_Cout, CIN 	=>	FA2_l5_c29_Cout, S =>	FA1_l4_c30_S, COUT 	=>	FA1_l4_c30_Cout );

	FA2_l4_c30  : FA 
	PORT MAP ( A =>	FA1_l5_c29_Cout, B =>	FA4_l5_c30_S, CIN 	=>	FA3_l5_c30_S, S =>	FA2_l4_c30_S, COUT 	=>	FA2_l4_c30_Cout );

	FA3_l4_c30  : FA 
	PORT MAP ( A =>	FA2_l5_c30_S, B =>	FA1_l5_c30_S, CIN 	=>	PP15(32), S =>	FA3_l4_c30_S, COUT 	=>	FA3_l4_c30_Cout );

	FA1_l4_c31  : FA
	PORT MAP ( A =>	FA4_l5_c30_Cout, B =>	FA3_l5_c30_Cout, CIN 	=>	FA2_l5_c30_Cout, S =>	FA1_l4_c31_S, COUT 	=>	FA1_l4_c31_Cout );

	FA2_l4_c31  : FA
	PORT MAP ( A =>	FA1_l5_c30_Cout, B =>	FA4_l5_c31_S, CIN 	=>	FA3_l5_c31_S, S =>	FA2_l4_c31_S, COUT 	=>	FA2_l4_c31_Cout );

	FA3_l4_c31  : FA 
	PORT MAP ( A =>	FA2_l5_c31_S, B =>	FA1_l5_c31_S, CIN 	=>	PP15(1), S =>	FA3_l4_c31_S, COUT 	=>	FA3_l4_c31_Cout );

	FA1_l4_c32  : FA 
	PORT MAP ( A =>	FA4_l5_c31_Cout, B =>	FA3_l5_c31_Cout, CIN 	=>	FA2_l5_c31_Cout, S =>	FA1_l4_c32_S, COUT 	=>	FA1_l4_c32_Cout );

	FA2_l4_c32  : FA 
	PORT MAP ( A =>	FA1_l5_c31_Cout, B =>	FA4_l5_c32_S, CIN 	=>	FA3_l5_c32_S, S =>	FA2_l4_c32_S, COUT 	=>	FA2_l4_c32_Cout );

	FA3_l4_c32  : FA 
	PORT MAP ( A =>	FA2_l5_c32_S, B =>	FA1_l5_c32_S, CIN 	=>	PP16(0), S =>	FA3_l4_c32_S, COUT 	=>	FA3_l4_c32_Cout );

	FA1_l4_c33  : FA 
	PORT MAP ( A =>	FA4_l5_c32_Cout, B =>	FA3_l5_c32_Cout, CIN 	=>	FA2_l5_c32_Cout, S =>	FA1_l4_c33_S, COUT 	=>	FA1_l4_c33_Cout );

	FA2_l4_c33  : FA 
	PORT MAP ( A =>	FA1_l5_c32_Cout, B =>	FA4_l5_c33_S, CIN 	=>	FA3_l5_c33_S, S =>	FA2_l4_c33_S, COUT 	=>	FA2_l4_c33_Cout );

	FA3_l4_c33  : FA 
	PORT MAP ( A =>	FA2_l5_c33_S, B =>	FA1_l5_c33_S, CIN 	=>	PP16(1), S =>	FA3_l4_c33_S, COUT 	=>	FA3_l4_c33_Cout );

	FA1_l4_c34  : FA 
	PORT MAP ( A =>	FA4_l5_c33_Cout, B =>	FA3_l5_c33_Cout, CIN 	=>	FA2_l5_c33_Cout, S =>	FA1_l4_c34_S, COUT 	=>	FA1_l4_c34_Cout );

	FA2_l4_c34  : FA 
	PORT MAP ( A =>	FA1_l5_c33_Cout, B =>	FA4_l5_c34_S, CIN 	=>	FA3_l5_c34_S, S =>	FA2_l4_c34_S, COUT 	=>	FA2_l4_c34_Cout );

	FA3_l4_c34  : FA 
	PORT MAP ( A =>	FA2_l5_c34_S, B =>	FA1_l5_c34_S, CIN 	=>	PP16(2), S =>	FA3_l4_c34_S, COUT 	=>	FA3_l4_c34_Cout );

	FA1_l4_c35  : FA 
	PORT MAP ( A =>	FA4_l5_c34_Cout, B =>	FA3_l5_c34_Cout, CIN 	=>	FA2_l5_c34_Cout, S =>	FA1_l4_c35_S, COUT 	=>	FA1_l4_c35_Cout );

	FA2_l4_c35  : FA 
	PORT MAP ( A =>	FA1_l5_c34_Cout, B =>	FA4_l5_c35_S, CIN 	=>	FA3_l5_c35_S, S =>	FA2_l4_c35_S, COUT 	=>	FA2_l4_c35_Cout );

	FA3_l4_c35  : FA 
	PORT MAP ( A =>	FA2_l5_c35_S, B =>	FA1_l5_c35_S, CIN 	=>	PP16(3), S =>	FA3_l4_c35_S, COUT 	=>	FA3_l4_c35_Cout );

	FA1_l4_c36  : FA 
	PORT MAP ( A =>	FA4_l5_c35_Cout, B =>	FA3_l5_c35_Cout, CIN 	=>	FA2_l5_c35_Cout, S =>	FA1_l4_c36_S, COUT 	=>	FA1_l4_c36_Cout );

	FA2_l4_c36  : FA 
	PORT MAP ( A =>	FA1_l5_c35_Cout, B =>	FA4_l5_c36_S, CIN 	=>	FA3_l5_c36_S, S =>	FA2_l4_c36_S, COUT 	=>	FA2_l4_c36_Cout );

	FA3_l4_c36  : FA 
	PORT MAP ( A =>	FA2_l5_c36_S, B =>	FA1_l5_c36_S, CIN 	=>	PP16(4), S =>	FA3_l4_c36_S, COUT 	=>	FA3_l4_c36_Cout );

	FA1_l4_c37  : FA 
	PORT MAP ( A =>	FA4_l5_c36_Cout, B =>	FA3_l5_c36_Cout, CIN 	=>	FA2_l5_c36_Cout, S =>	FA1_l4_c37_S, COUT 	=>	FA1_l4_c37_Cout );

	FA2_l4_c37  : FA 
	PORT MAP ( A =>	FA1_l5_c36_Cout, B =>	FA4_l5_c37_S, CIN 	=>	FA3_l5_c37_S, S =>	FA2_l4_c37_S, COUT 	=>	FA2_l4_c37_Cout );

	FA3_l4_c37  : FA 
	PORT MAP ( A =>	FA2_l5_c37_S, B =>	FA1_l5_c37_S, CIN 	=>	PP16(5), S =>	FA3_l4_c37_S, COUT 	=>	FA3_l4_c37_Cout );

	FA1_l4_c38  : FA 
	PORT MAP ( A =>	FA4_l5_c37_Cout, B =>	FA3_l5_c37_Cout, CIN 	=>	FA2_l5_c37_Cout, S =>	FA1_l4_c38_S, COUT 	=>	FA1_l4_c38_Cout );

	FA2_l4_c38  : FA 
	PORT MAP ( A =>	FA1_l5_c37_Cout, B =>	FA4_l5_c38_S, CIN 	=>	FA3_l5_c38_S, S =>	FA2_l4_c38_S, COUT 	=>	FA2_l4_c38_Cout );

	FA3_l4_c38  : FA 
	PORT MAP ( A =>	FA2_l5_c38_S, B =>	FA1_l5_c38_S, CIN 	=>	PP16(6), S =>	FA3_l4_c38_S, COUT 	=>	FA3_l4_c38_Cout );

	FA1_l4_c39  : FA 
	PORT MAP ( A =>	FA4_l5_c38_Cout, B =>	FA3_l5_c38_Cout, CIN 	=>	FA2_l5_c38_Cout, S =>	FA1_l4_c39_S, COUT 	=>	FA1_l4_c39_Cout );

	FA2_l4_c39  : FA 
	PORT MAP ( A =>	FA1_l5_c38_Cout, B =>	FA4_l5_c39_S, CIN 	=>	FA3_l5_c39_S, S =>	FA2_l4_c39_S, COUT 	=>	FA2_l4_c39_Cout );

	FA3_l4_c39  : FA 
	PORT MAP ( A =>	FA2_l5_c39_S, B =>	FA1_l5_c39_S, CIN 	=>	PP16(7), S =>	FA3_l4_c39_S, COUT 	=>	FA3_l4_c39_Cout );

	FA1_l4_c40  : FA 
	PORT MAP ( A =>	FA4_l5_c39_Cout, B =>	FA3_l5_c39_Cout, CIN 	=>	FA2_l5_c39_Cout, S =>	FA1_l4_c40_S, COUT 	=>	FA1_l4_c40_Cout );

	FA2_l4_c40  : FA 
	PORT MAP ( A =>	FA1_l5_c39_Cout, B =>	FA4_l5_c40_S, CIN 	=>	FA3_l5_c40_S, S =>	FA2_l4_c40_S, COUT 	=>	FA2_l4_c40_Cout );

	FA3_l4_c40  : FA 
	PORT MAP ( A =>	FA2_l5_c40_S, B =>	FA1_l5_c40_S, CIN 	=>	PP16(8), S =>	FA3_l4_c40_S, COUT 	=>	FA3_l4_c40_Cout );

	FA1_l4_c41  : FA 
	PORT MAP ( A =>	FA4_l5_c40_Cout, B =>	FA3_l5_c40_Cout, CIN 	=>	FA2_l5_c40_Cout, S =>	FA1_l4_c41_S, COUT 	=>	FA1_l4_c41_Cout );

	FA2_l4_c41  : FA 
	PORT MAP ( A =>	FA1_l5_c40_Cout, B =>	FA4_l5_c41_S, CIN 	=>	FA3_l5_c41_S, S =>	FA2_l4_c41_S, COUT 	=>	FA2_l4_c41_Cout );

	FA3_l4_c41  : FA 
	PORT MAP ( A =>	FA2_l5_c41_S, B =>	FA1_l5_c41_S, CIN 	=>	PP16(9), S =>	FA3_l4_c41_S, COUT 	=>	FA3_l4_c41_Cout );

	FA1_l4_c42  : FA 
	PORT MAP ( A =>	FA4_l5_c41_Cout, B =>	FA3_l5_c41_Cout, CIN 	=>	FA2_l5_c41_Cout, S =>	FA1_l4_c42_S, COUT 	=>	FA1_l4_c42_Cout );

	FA2_l4_c42  : FA 
	PORT MAP ( A =>	FA1_l5_c41_Cout, B =>	FA4_l5_c42_S, CIN 	=>	FA3_l5_c42_S, S =>	FA2_l4_c42_S, COUT 	=>	FA2_l4_c42_Cout );

	FA3_l4_c42  : FA
	PORT MAP ( A =>	FA2_l5_c42_S, B =>	FA1_l5_c42_S, CIN 	=>	PP16(10), S =>	FA3_l4_c42_S, COUT 	=>	FA3_l4_c42_Cout );

	FA1_l4_c43  : FA 
	PORT MAP ( A =>	FA4_l5_c42_Cout, B =>	FA3_l5_c42_Cout, CIN 	=>	FA2_l5_c42_Cout, S =>	FA1_l4_c43_S, COUT 	=>	FA1_l4_c43_Cout );

	FA2_l4_c43  : FA 
	PORT MAP ( A =>	FA1_l5_c42_Cout, B =>	FA4_l5_c43_S, CIN 	=>	FA3_l5_c43_S, S =>	FA2_l4_c43_S, COUT 	=>	FA2_l4_c43_Cout );

	FA3_l4_c43  : FA 
	PORT MAP ( A =>	FA2_l5_c43_S, B =>	FA1_l5_c43_S, CIN 	=>	PP16(11), S =>	FA3_l4_c43_S, COUT 	=>	FA3_l4_c43_Cout );

	FA1_l4_c44  : FA 
	PORT MAP ( A =>	FA4_l5_c43_Cout, B =>	FA3_l5_c43_Cout, CIN 	=>	FA2_l5_c43_Cout, S =>	FA1_l4_c44_S, COUT 	=>	FA1_l4_c44_Cout );

	FA2_l4_c44  : FA 
	PORT MAP ( A =>	FA1_l5_c43_Cout, B =>	HA1_l5_c44_S, CIN 	=>	FA3_l5_c44_S, S =>	FA2_l4_c44_S, COUT 	=>	FA2_l4_c44_Cout );

	FA3_l4_c44  : FA 
	PORT MAP ( A =>	FA2_l5_c44_S, B =>	FA1_l5_c44_S, CIN 	=>	PP16(12), S =>	FA3_l4_c44_S, COUT 	=>	FA3_l4_c44_Cout );

	FA1_l4_c45  : FA 
	PORT MAP ( A =>	HA1_l5_c44_Cout, B =>	FA3_l5_c44_Cout, CIN 	=>	FA2_l5_c44_Cout, S =>	FA1_l4_c45_S, COUT 	=>	FA1_l4_c45_Cout );

	FA2_l4_c45  : FA 
	PORT MAP ( A =>	FA1_l5_c44_Cout, B =>	FA3_l5_c45_S, CIN 	=>	FA2_l5_c45_S, S =>	FA2_l4_c45_S, COUT 	=>	FA2_l4_c45_Cout );

	FA3_l4_c45  : FA 
	PORT MAP ( A =>	FA1_l5_c45_S, B =>	PP15(15), CIN 	=>	PP16(13), S =>	FA3_l4_c45_S, COUT 	=>	FA3_l4_c45_Cout );

	FA1_l4_c46  : FA 
	PORT MAP ( A =>	FA3_l5_c45_Cout, B =>	FA2_l5_c45_Cout, CIN 	=>	FA1_l5_c45_Cout, S =>	FA1_l4_c46_S, COUT 	=>	FA1_l4_c46_Cout );

	FA2_l4_c46  : FA 
	PORT MAP ( A =>	HA1_l5_c46_S, B =>	FA2_l5_c46_S, CIN 	=>	FA1_l5_c46_S, S =>	FA2_l4_c46_S, COUT 	=>	FA2_l4_c46_Cout );

	FA3_l4_c46  : FA 
	PORT MAP ( A =>	PP14(18), B =>	PP15(16), CIN 	=>	PP16(14), S =>	FA3_l4_c46_S, COUT 	=>	FA3_l4_c46_Cout );

	FA1_l4_c47  : FA 
	PORT MAP ( A =>	HA1_l5_c46_Cout, B =>	FA2_l5_c46_Cout, CIN 	=>	FA1_l5_c46_Cout, S =>	FA1_l4_c47_S, COUT 	=>	FA1_l4_c47_Cout );

	FA2_l4_c47  : FA 
	PORT MAP ( A =>	FA2_l5_c47_S, B =>	FA1_l5_c47_S, CIN 	=>	PP13(21), S =>	FA2_l4_c47_S, COUT 	=>	FA2_l4_c47_Cout );

	FA3_l4_c47  : FA 
	PORT MAP ( A =>	PP14(19), B =>	PP15(17), CIN 	=>	PP16(15), S =>	FA3_l4_c47_S, COUT 	=>	FA3_l4_c47_Cout );

	FA1_l4_c48  : FA 
	PORT MAP ( A =>	FA2_l5_c47_Cout, B =>	FA1_l5_c47_Cout, CIN 	=>	HA1_l5_c48_S, S =>	FA1_l4_c48_S, COUT 	=>	FA1_l4_c48_Cout );

	FA2_l4_c48  : FA 
	PORT MAP ( A =>	FA1_l5_c48_S, B =>	PP12(24), CIN 	=>	PP13(22), S =>	FA2_l4_c48_S, COUT 	=>	FA2_l4_c48_Cout );

	FA3_l4_c48  : FA 
	PORT MAP ( A =>	PP14(20), B =>	PP15(18), CIN 	=>	PP16(16), S =>	FA3_l4_c48_S, COUT 	=>	FA3_l4_c48_Cout );

	FA1_l4_c49  : FA 
	PORT MAP ( A =>	HA1_l5_c48_Cout, B =>	FA1_l5_c48_Cout, CIN 	=>	FA1_l5_c49_S, S =>	FA1_l4_c49_S, COUT 	=>	FA1_l4_c49_Cout );

	FA2_l4_c49  : FA 
	PORT MAP ( A =>	PP11(27), B =>	PP12(25), CIN 	=>	PP13(23), S =>	FA2_l4_c49_S, COUT 	=>	FA2_l4_c49_Cout );

	FA3_l4_c49  : FA 
	PORT MAP ( A =>	PP14(21), B =>	PP15(19), CIN 	=>	PP16(17), S =>	FA3_l4_c49_S, COUT 	=>	FA3_l4_c49_Cout );

	FA1_l4_c50  : FA 
	PORT MAP ( A =>	FA1_l5_c49_Cout, B =>	HA1_l5_c50_S, CIN 	=>	PP10(30), S =>	FA1_l4_c50_S, COUT 	=>	FA1_l4_c50_Cout );

	FA2_l4_c50  : FA 
	PORT MAP ( A =>	PP11(28), B =>	PP12(26), CIN 	=>	PP13(24), S =>	FA2_l4_c50_S, COUT 	=>	FA2_l4_c50_Cout );

	FA3_l4_c50  : FA 
	PORT MAP ( A =>	PP14(22), B =>	PP15(20), CIN 	=>	PP16(18), S =>	FA3_l4_c50_S, COUT 	=>	FA3_l4_c50_Cout );

	FA1_l4_c51  : FA 
	PORT MAP ( A =>	HA1_l5_c50_Cout, B =>	PP9_neg, CIN 	=>	PP10(31), S =>	FA1_l4_c51_S, COUT 	=>	FA1_l4_c51_Cout );

	FA2_l4_c51  : FA 
	PORT MAP ( A =>	PP11(29), B =>	PP12(27), CIN 	=>	PP13(25), S =>	FA2_l4_c51_S, COUT 	=>	FA2_l4_c51_Cout );

	FA3_l4_c51  : FA 
	PORT MAP ( A =>	PP14(23), B =>	PP15(21), CIN 	=>	PP16(19), S =>	FA3_l4_c51_S, COUT 	=>	FA3_l4_c51_Cout );

	FA1_l4_c52  : FA
	PORT MAP ( A =>	'1', B =>	PP10(32), CIN 	=>	PP11(30), S =>	FA1_l4_c52_S, COUT 	=>	FA1_l4_c52_Cout );

	FA2_l4_c52  : FA 
	PORT MAP ( A =>	PP12(28), B =>	PP13(26), CIN 	=>	PP14(24), S =>	FA2_l4_c52_S, COUT 	=>	FA2_l4_c52_Cout );

	HA1_l4_c52  : HA 
	PORT MAP ( A =>	PP15(22), B =>	PP16(20), S =>	HA1_l4_c52_S, COUT 	=>	HA1_l4_c52_Cout );

	FA1_l4_c53  : FA 
	PORT MAP ( A =>	PP10_neg, B =>	PP11(31), CIN 	=>	PP12(29), S =>	FA1_l4_c53_S, COUT 	=>	FA1_l4_c53_Cout );

	FA2_l4_c53  : FA 
	PORT MAP ( A =>	PP13(27), B =>	PP14(25), CIN 	=>	PP15(23), S =>	FA2_l4_c53_S, COUT 	=>	FA2_l4_c53_Cout );

	FA1_l4_c54  : FA 
	PORT MAP ( A =>	'1', B =>	PP11(32), CIN 	=>	PP12(30), S =>	FA1_l4_c54_S, COUT 	=>	FA1_l4_c54_Cout );

	HA1_l4_c54  : HA 
	PORT MAP ( A =>	PP13(28), B =>	PP14(26), S =>	HA1_l4_c54_S, COUT 	=>	HA1_l4_c54_Cout );

	FA1_l4_c55  : FA 
	PORT MAP ( A =>	PP11_neg, B =>	PP12(31), CIN 	=>	PP13(29), S =>	FA1_l4_c55_S, COUT 	=>	FA1_l4_c55_Cout );

	HA1_l4_c56  : HA 
	PORT MAP ( A =>	'1', B =>	PP12(32), S =>	HA1_l4_c56_S, COUT 	=>	HA1_l4_c56_Cout );

	HA1_l3_c6  : HA 
	PORT MAP ( A =>	PP0(6), B =>	PP1(4), S =>	HA1_l3_c6_S, COUT 	=>	HA1_l3_c6_Cout );

	HA1_l3_c7  : HA 
	PORT MAP ( A =>	PP0(7), B =>	PP1(5), S =>	HA1_l3_c7_S, COUT 	=>	HA1_l3_c7_Cout );

	FA1_l3_c8  : FA 
	PORT MAP ( A =>	PP0(8), B =>	PP1(6), CIN 	=>	PP2(4), S =>	FA1_l3_c8_S, COUT 	=>	FA1_l3_c8_Cout );

	HA1_l3_c8  : HA 
	PORT MAP ( A =>	PP3(2), B =>	PP4(0), S =>	HA1_l3_c8_S, COUT 	=>	HA1_l3_c8_Cout );

	FA1_l3_c9  : FA 
	PORT MAP ( A =>	PP0(9), B =>	PP1(7), CIN 	=>	PP2(5), S =>	FA1_l3_c9_S, COUT 	=>	FA1_l3_c9_Cout );

	HA1_l3_c9  : HA 
	PORT MAP ( A =>	PP3(3), B =>	PP4(1), S =>	HA1_l3_c9_S, COUT 	=>	HA1_l3_c9_Cout );

	FA1_l3_c10  : FA 
	PORT MAP ( A =>	HA1_l4_c10_S, B =>	PP2(6), CIN 	=>	PP3(4), S =>	FA1_l3_c10_S, COUT 	=>	FA1_l3_c10_Cout );

	FA2_l3_c10  : FA
	PORT MAP ( A =>	PP4(2), B =>	PP5(0), CIN 	=>	PP5(32), S =>	FA2_l3_c10_S, COUT 	=>	FA2_l3_c10_Cout );

	FA1_l3_c11  : FA 
	PORT MAP ( A =>	HA1_l4_c10_Cout, B =>	HA1_l4_c11_S, CIN 	=>	PP2(7), S =>	FA1_l3_c11_S, COUT 	=>	FA1_l3_c11_Cout );

	FA2_l3_c11  : FA 
	PORT MAP ( A =>	PP3(5), B =>	PP4(3), CIN 	=>	PP5(1), S =>	FA2_l3_c11_S, COUT 	=>	FA2_l3_c11_Cout );

	FA1_l3_c12  : FA 
	PORT MAP ( A =>	HA1_l4_c11_Cout, B =>	HA1_l4_c12_S, CIN 	=>	FA1_l4_c12_S, S =>	FA1_l3_c12_S, COUT 	=>	FA1_l3_c12_Cout );

	FA2_l3_c12  : FA 
	PORT MAP ( A =>	PP5(2), B =>	PP6(0), CIN 	=>	PP6(32), S =>	FA2_l3_c12_S, COUT 	=>	FA2_l3_c12_Cout );

	FA1_l3_c13  : FA 
	PORT MAP ( A =>	HA1_l4_c12_Cout, B =>	FA1_l4_c12_Cout, CIN 	=>	HA1_l4_c13_S, S =>	FA1_l3_c13_S, COUT 	=>	FA1_l3_c13_Cout );

	FA2_l3_c13  : FA 
	PORT MAP ( A =>	FA1_l4_c13_S, B =>	PP5(3), CIN 	=>	PP6(1), S =>	FA2_l3_c13_S, COUT 	=>	FA2_l3_c13_Cout );

	FA1_l3_c14  : FA 
	PORT MAP ( A =>	HA1_l4_c13_Cout, B =>	FA1_l4_c13_Cout, CIN 	=>	HA1_l4_c14_S, S =>	FA1_l3_c14_S, COUT 	=>	FA1_l3_c14_Cout );

	FA2_l3_c14  : FA 
	PORT MAP ( A =>	FA2_l4_c14_S, B =>	FA1_l4_c14_S, CIN 	=>	PP7(32), S =>	FA2_l3_c14_S, COUT 	=>	FA2_l3_c14_Cout );

	FA1_l3_c15  : FA 
	PORT MAP ( A =>	HA1_l4_c14_Cout, B =>	FA2_l4_c14_Cout, CIN 	=>	FA1_l4_c14_Cout, S =>	FA1_l3_c15_S, COUT 	=>	FA1_l3_c15_Cout );

	FA2_l3_c15  : FA 
	PORT MAP ( A =>	HA1_l4_c15_S, B =>	FA2_l4_c15_S, CIN 	=>	FA1_l4_c15_S, S =>	FA2_l3_c15_S, COUT 	=>	FA2_l3_c15_Cout );

	FA1_l3_c16  : FA 
	PORT MAP ( A =>	HA1_l4_c15_Cout, B =>	FA2_l4_c15_Cout, CIN 	=>	FA1_l4_c15_Cout, S =>	FA1_l3_c16_S, COUT 	=>	FA1_l3_c16_Cout );

	FA2_l3_c16  : FA
	PORT MAP ( A =>	FA3_l4_c16_S, B =>	FA2_l4_c16_S, CIN 	=>	FA1_l4_c16_S, S =>	FA2_l3_c16_S, COUT 	=>	FA2_l3_c16_Cout );

	FA1_l3_c17  : FA 
	PORT MAP ( A =>	FA3_l4_c16_Cout, B =>	FA2_l4_c16_Cout, CIN 	=>	FA1_l4_c16_Cout, S =>	FA1_l3_c17_S, COUT 	=>	FA1_l3_c17_Cout );

	FA2_l3_c17  : FA 
	PORT MAP ( A =>	FA3_l4_c17_S, B =>	FA2_l4_c17_S, CIN 	=>	FA1_l4_c17_S, S =>	FA2_l3_c17_S, COUT 	=>	FA2_l3_c17_Cout );

	FA1_l3_c18  : FA 
	PORT MAP ( A =>	FA3_l4_c17_Cout, B =>	FA2_l4_c17_Cout, CIN 	=>	FA1_l4_c17_Cout, S =>	FA1_l3_c18_S, COUT 	=>	FA1_l3_c18_Cout );

	FA2_l3_c18  : FA 
	PORT MAP ( A =>	FA3_l4_c18_S, B =>	FA2_l4_c18_S, CIN 	=>	FA1_l4_c18_S, S =>	FA2_l3_c18_S, COUT 	=>	FA2_l3_c18_Cout );

	FA1_l3_c19  : FA 
	PORT MAP ( A =>	FA3_l4_c18_Cout, B =>	FA2_l4_c18_Cout, CIN 	=>	FA1_l4_c18_Cout, S =>	FA1_l3_c19_S, COUT 	=>	FA1_l3_c19_Cout );

	FA2_l3_c19  : FA 
	PORT MAP ( A =>	FA3_l4_c19_S, B =>	FA2_l4_c19_S, CIN 	=>	FA1_l4_c19_S, S =>	FA2_l3_c19_S, COUT 	=>	FA2_l3_c19_Cout );

	FA1_l3_c20  : FA 
	PORT MAP ( A =>	FA3_l4_c19_Cout, B =>	FA2_l4_c19_Cout, CIN 	=>	FA1_l4_c19_Cout, S =>	FA1_l3_c20_S, COUT 	=>	FA1_l3_c20_Cout );

	FA2_l3_c20  : FA 
	PORT MAP ( A =>	FA3_l4_c20_S, B =>	FA2_l4_c20_S, CIN 	=>	FA1_l4_c20_S, S =>	FA2_l3_c20_S, COUT 	=>	FA2_l3_c20_Cout );

	FA1_l3_c21  : FA 
	PORT MAP ( A =>	FA3_l4_c20_Cout, B =>	FA2_l4_c20_Cout, CIN 	=>	FA1_l4_c20_Cout, S =>	FA1_l3_c21_S, COUT 	=>	FA1_l3_c21_Cout );

	FA2_l3_c21  : FA 
	PORT MAP ( A =>	FA3_l4_c21_S, B =>	FA2_l4_c21_S, CIN 	=>	FA1_l4_c21_S, S =>	FA2_l3_c21_S, COUT 	=>	FA2_l3_c21_Cout );

	FA1_l3_c22  : FA 
	PORT MAP ( A =>	FA3_l4_c21_Cout, B =>	FA2_l4_c21_Cout, CIN 	=>	FA1_l4_c21_Cout, S =>	FA1_l3_c22_S, COUT 	=>	FA1_l3_c22_Cout );

	FA2_l3_c22  : FA 
	PORT MAP ( A =>	FA3_l4_c22_S, B =>	FA2_l4_c22_S, CIN 	=>	FA1_l4_c22_S, S =>	FA2_l3_c22_S, COUT 	=>	FA2_l3_c22_Cout );

	FA1_l3_c23  : FA 
	PORT MAP ( A =>	FA3_l4_c22_Cout, B =>	FA2_l4_c22_Cout, CIN 	=>	FA1_l4_c22_Cout, S =>	FA1_l3_c23_S, COUT 	=>	FA1_l3_c23_Cout );

	FA2_l3_c23  : FA 
	PORT MAP ( A =>	FA3_l4_c23_S, B =>	FA2_l4_c23_S, CIN 	=>	FA1_l4_c23_S, S =>	FA2_l3_c23_S, COUT 	=>	FA2_l3_c23_Cout );

	FA1_l3_c24  : FA 
	PORT MAP ( A =>	FA3_l4_c23_Cout, B =>	FA2_l4_c23_Cout, CIN 	=>	FA1_l4_c23_Cout, S =>	FA1_l3_c24_S, COUT 	=>	FA1_l3_c24_Cout );

	FA2_l3_c24  : FA 
	PORT MAP ( A =>	FA3_l4_c24_S, B =>	FA2_l4_c24_S, CIN 	=>	FA1_l4_c24_S, S =>	FA2_l3_c24_S, COUT 	=>	FA2_l3_c24_Cout );

	FA1_l3_c25  : FA 
	PORT MAP ( A =>	FA3_l4_c24_Cout, B =>	FA2_l4_c24_Cout, CIN 	=>	FA1_l4_c24_Cout, S =>	FA1_l3_c25_S, COUT 	=>	FA1_l3_c25_Cout );

	FA2_l3_c25  : FA 
	PORT MAP ( A =>	FA3_l4_c25_S, B =>	FA2_l4_c25_S, CIN 	=>	FA1_l4_c25_S, S =>	FA2_l3_c25_S, COUT 	=>	FA2_l3_c25_Cout );

	FA1_l3_c26  : FA 
	PORT MAP ( A =>	FA3_l4_c25_Cout, B =>	FA2_l4_c25_Cout, CIN 	=>	FA1_l4_c25_Cout, S =>	FA1_l3_c26_S, COUT 	=>	FA1_l3_c26_Cout );

	FA2_l3_c26  : FA 
	PORT MAP ( A =>	FA3_l4_c26_S, B =>	FA2_l4_c26_S, CIN 	=>	FA1_l4_c26_S, S =>	FA2_l3_c26_S, COUT 	=>	FA2_l3_c26_Cout );

	FA1_l3_c27  : FA 
	PORT MAP ( A =>	FA3_l4_c26_Cout, B =>	FA2_l4_c26_Cout, CIN 	=>	FA1_l4_c26_Cout, S =>	FA1_l3_c27_S, COUT 	=>	FA1_l3_c27_Cout );

	FA2_l3_c27  : FA 
	PORT MAP ( A =>	FA3_l4_c27_S, B =>	FA2_l4_c27_S, CIN 	=>	FA1_l4_c27_S, S =>	FA2_l3_c27_S, COUT 	=>	FA2_l3_c27_Cout );

	FA1_l3_c28  : FA 
	PORT MAP ( A =>	FA3_l4_c27_Cout, B =>	FA2_l4_c27_Cout, CIN 	=>	FA1_l4_c27_Cout, S =>	FA1_l3_c28_S, COUT 	=>	FA1_l3_c28_Cout );

	FA2_l3_c28  : FA 
	PORT MAP ( A =>	FA3_l4_c28_S, B =>	FA2_l4_c28_S, CIN 	=>	FA1_l4_c28_S, S =>	FA2_l3_c28_S, COUT 	=>	FA2_l3_c28_Cout );

	FA1_l3_c29  : FA 
	PORT MAP ( A =>	FA3_l4_c28_Cout, B =>	FA2_l4_c28_Cout, CIN 	=>	FA1_l4_c28_Cout, S =>	FA1_l3_c29_S, COUT 	=>	FA1_l3_c29_Cout );

	FA2_l3_c29  : FA 
	PORT MAP ( A =>	FA3_l4_c29_S, B =>	FA2_l4_c29_S, CIN 	=>	FA1_l4_c29_S, S =>	FA2_l3_c29_S, COUT 	=>	FA2_l3_c29_Cout );

	FA1_l3_c30  : FA 
	PORT MAP ( A =>	FA3_l4_c29_Cout, B =>	FA2_l4_c29_Cout, CIN 	=>	FA1_l4_c29_Cout, S =>	FA1_l3_c30_S, COUT 	=>	FA1_l3_c30_Cout );

	FA2_l3_c30  : FA 
	PORT MAP ( A =>	FA3_l4_c30_S, B =>	FA2_l4_c30_S, CIN 	=>	FA1_l4_c30_S, S =>	FA2_l3_c30_S, COUT 	=>	FA2_l3_c30_Cout );

	FA1_l3_c31  : FA 
	PORT MAP ( A =>	FA3_l4_c30_Cout, B =>	FA2_l4_c30_Cout, CIN 	=>	FA1_l4_c30_Cout, S =>	FA1_l3_c31_S, COUT 	=>	FA1_l3_c31_Cout );

	FA2_l3_c31  : FA 
	PORT MAP ( A =>	FA3_l4_c31_S, B =>	FA2_l4_c31_S, CIN 	=>	FA1_l4_c31_S, S =>	FA2_l3_c31_S, COUT 	=>	FA2_l3_c31_Cout );

	FA1_l3_c32  : FA 
	PORT MAP ( A =>	FA3_l4_c31_Cout, B =>	FA2_l4_c31_Cout, CIN 	=>	FA1_l4_c31_Cout, S =>	FA1_l3_c32_S, COUT 	=>	FA1_l3_c32_Cout );

	FA2_l3_c32  : FA 
	PORT MAP ( A =>	FA3_l4_c32_S, B =>	FA2_l4_c32_S, CIN 	=>	FA1_l4_c32_S, S =>	FA2_l3_c32_S, COUT 	=>	FA2_l3_c32_Cout );

	FA1_l3_c33  : FA
	PORT MAP ( A =>	FA3_l4_c32_Cout, B =>	FA2_l4_c32_Cout, CIN 	=>	FA1_l4_c32_Cout, S =>	FA1_l3_c33_S, COUT 	=>	FA1_l3_c33_Cout );

	FA2_l3_c33  : FA 
	PORT MAP ( A =>	FA3_l4_c33_S, B =>	FA2_l4_c33_S, CIN 	=>	FA1_l4_c33_S, S =>	FA2_l3_c33_S, COUT 	=>	FA2_l3_c33_Cout );

	FA1_l3_c34  : FA 
	PORT MAP ( A =>	FA3_l4_c33_Cout, B =>	FA2_l4_c33_Cout, CIN 	=>	FA1_l4_c33_Cout, S =>	FA1_l3_c34_S, COUT 	=>	FA1_l3_c34_Cout );
	
	FA2_l3_c34  : FA 
	PORT MAP ( A =>	FA3_l4_c34_S, B =>	FA2_l4_c34_S, CIN 	=>	FA1_l4_c34_S, S =>	FA2_l3_c34_S, COUT 	=>	FA2_l3_c34_Cout );

	FA1_l3_c35  : FA 
	PORT MAP ( A =>	FA3_l4_c34_Cout, B =>	FA2_l4_c34_Cout, CIN 	=>	FA1_l4_c34_Cout, S =>	FA1_l3_c35_S, COUT 	=>	FA1_l3_c35_Cout );

	FA2_l3_c35  : FA 
	PORT MAP ( A =>	FA3_l4_c35_S, B =>	FA2_l4_c35_S, CIN 	=>	FA1_l4_c35_S, S =>	FA2_l3_c35_S, COUT 	=>	FA2_l3_c35_Cout );

	FA1_l3_c36  : FA
	PORT MAP ( A =>	FA3_l4_c35_Cout, B =>	FA2_l4_c35_Cout, CIN 	=>	FA1_l4_c35_Cout, S =>	FA1_l3_c36_S, COUT 	=>	FA1_l3_c36_Cout );

	FA2_l3_c36  : FA 
	PORT MAP ( A =>	FA3_l4_c36_S, B =>	FA2_l4_c36_S, CIN 	=>	FA1_l4_c36_S, S =>	FA2_l3_c36_S, COUT 	=>	FA2_l3_c36_Cout );

	FA1_l3_c37  : FA 
	PORT MAP ( A =>	FA3_l4_c36_Cout, B =>	FA2_l4_c36_Cout, CIN 	=>	FA1_l4_c36_Cout, S =>	FA1_l3_c37_S, COUT 	=>	FA1_l3_c37_Cout );

	FA2_l3_c37  : FA
	PORT MAP ( A =>	FA3_l4_c37_S, B =>	FA2_l4_c37_S, CIN 	=>	FA1_l4_c37_S, S =>	FA2_l3_c37_S, COUT 	=>	FA2_l3_c37_Cout );

	FA1_l3_c38  : FA 
	PORT MAP ( A =>	FA3_l4_c37_Cout, B =>	FA2_l4_c37_Cout, CIN 	=>	FA1_l4_c37_Cout, S =>	FA1_l3_c38_S, COUT 	=>	FA1_l3_c38_Cout );

	FA2_l3_c38  : FA 
	PORT MAP ( A =>	FA3_l4_c38_S, B =>	FA2_l4_c38_S, CIN 	=>	FA1_l4_c38_S, S =>	FA2_l3_c38_S, COUT 	=>	FA2_l3_c38_Cout );

	FA1_l3_c39  : FA
	PORT MAP ( A =>	FA3_l4_c38_Cout, B =>	FA2_l4_c38_Cout, CIN 	=>	FA1_l4_c38_Cout, S =>	FA1_l3_c39_S, COUT 	=>	FA1_l3_c39_Cout );

	FA2_l3_c39  : FA
	PORT MAP ( A =>	FA3_l4_c39_S, B =>	FA2_l4_c39_S, CIN 	=>	FA1_l4_c39_S, S =>	FA2_l3_c39_S, COUT 	=>	FA2_l3_c39_Cout );

	FA1_l3_c40  : FA 
	PORT MAP ( A =>	FA3_l4_c39_Cout, B =>	FA2_l4_c39_Cout, CIN 	=>	FA1_l4_c39_Cout, S =>	FA1_l3_c40_S, COUT 	=>	FA1_l3_c40_Cout );

	FA2_l3_c40  : FA 
	PORT MAP ( A =>	FA3_l4_c40_S, B =>	FA2_l4_c40_S, CIN 	=>	FA1_l4_c40_S, S =>	FA2_l3_c40_S, COUT 	=>	FA2_l3_c40_Cout );

	FA1_l3_c41  : FA 
	PORT MAP ( A =>	FA3_l4_c40_Cout, B =>	FA2_l4_c40_Cout, CIN 	=>	FA1_l4_c40_Cout, S =>	FA1_l3_c41_S, COUT 	=>	FA1_l3_c41_Cout );

	FA2_l3_c41  : FA 
	PORT MAP ( A =>	FA3_l4_c41_S, B =>	FA2_l4_c41_S, CIN 	=>	FA1_l4_c41_S, S =>	FA2_l3_c41_S, COUT 	=>	FA2_l3_c41_Cout );

	FA1_l3_c42  : FA 
	PORT MAP ( A =>	FA3_l4_c41_Cout, B =>	FA2_l4_c41_Cout, CIN 	=>	FA1_l4_c41_Cout, S =>	FA1_l3_c42_S, COUT 	=>	FA1_l3_c42_Cout );

	FA2_l3_c42  : FA 
	PORT MAP ( A =>	FA3_l4_c42_S, B =>	FA2_l4_c42_S, CIN 	=>	FA1_l4_c42_S, S =>	FA2_l3_c42_S, COUT 	=>	FA2_l3_c42_Cout );

	FA1_l3_c43  : FA 
	PORT MAP ( A =>	FA3_l4_c42_Cout, B =>	FA2_l4_c42_Cout, CIN 	=>	FA1_l4_c42_Cout, S =>	FA1_l3_c43_S, COUT 	=>	FA1_l3_c43_Cout );

	FA2_l3_c43  : FA 
	PORT MAP ( A =>	FA3_l4_c43_S, B =>	FA2_l4_c43_S, CIN 	=>	FA1_l4_c43_S, S =>	FA2_l3_c43_S, COUT 	=>	FA2_l3_c43_Cout );

	FA1_l3_c44  : FA 
	PORT MAP ( A =>	FA3_l4_c43_Cout, B =>	FA2_l4_c43_Cout, CIN 	=>	FA1_l4_c43_Cout, S =>	FA1_l3_c44_S, COUT 	=>	FA1_l3_c44_Cout );

	FA2_l3_c44  : FA 
	PORT MAP ( A =>	FA3_l4_c44_S, B =>	FA2_l4_c44_S, CIN 	=>	FA1_l4_c44_S, S =>	FA2_l3_c44_S, COUT 	=>	FA2_l3_c44_Cout );

	FA1_l3_c45  : FA 
	PORT MAP ( A =>	FA3_l4_c44_Cout, B =>	FA2_l4_c44_Cout, CIN 	=>	FA1_l4_c44_Cout, S =>	FA1_l3_c45_S, COUT 	=>	FA1_l3_c45_Cout );

	FA2_l3_c45  : FA 
	PORT MAP ( A =>	FA3_l4_c45_S, B =>	FA2_l4_c45_S, CIN 	=>	FA1_l4_c45_S, S =>	FA2_l3_c45_S, COUT 	=>	FA2_l3_c45_Cout );

	FA1_l3_c46  : FA 
	PORT MAP ( A =>	FA3_l4_c45_Cout, B =>	FA2_l4_c45_Cout, CIN 	=>	FA1_l4_c45_Cout, S =>	FA1_l3_c46_S, COUT 	=>	FA1_l3_c46_Cout );

	FA2_l3_c46  : FA 
	PORT MAP ( A =>	FA3_l4_c46_S, B =>	FA2_l4_c46_S, CIN 	=>	FA1_l4_c46_S, S =>	FA2_l3_c46_S, COUT 	=>	FA2_l3_c46_Cout );

	FA1_l3_c47  : FA 
	PORT MAP ( A =>	FA3_l4_c46_Cout, B =>	FA2_l4_c46_Cout, CIN 	=>	FA1_l4_c46_Cout, S =>	FA1_l3_c47_S, COUT 	=>	FA1_l3_c47_Cout );

	FA2_l3_c47  : FA 
	PORT MAP ( A =>	FA3_l4_c47_S, B =>	FA2_l4_c47_S, CIN 	=>	FA1_l4_c47_S, S =>	FA2_l3_c47_S, COUT 	=>	FA2_l3_c47_Cout );

	FA1_l3_c48  : FA 
	PORT MAP ( A =>	FA3_l4_c47_Cout, B =>	FA2_l4_c47_Cout, CIN 	=>	FA1_l4_c47_Cout, S =>	FA1_l3_c48_S, COUT 	=>	FA1_l3_c48_Cout );

	FA2_l3_c48  : FA 
	PORT MAP ( A =>	FA3_l4_c48_S, B =>	FA2_l4_c48_S, CIN 	=>	FA1_l4_c48_S, S =>	FA2_l3_c48_S, COUT 	=>	FA2_l3_c48_Cout );

	FA1_l3_c49  : FA 
	PORT MAP ( A =>	FA3_l4_c48_Cout, B =>	FA2_l4_c48_Cout, CIN 	=>	FA1_l4_c48_Cout, S =>	FA1_l3_c49_S, COUT 	=>	FA1_l3_c49_Cout );

	FA2_l3_c49  : FA 
	PORT MAP ( A =>	FA3_l4_c49_S, B =>	FA2_l4_c49_S, CIN 	=>	FA1_l4_c49_S, S =>	FA2_l3_c49_S, COUT 	=>	FA2_l3_c49_Cout );

	FA1_l3_c50  : FA 
	PORT MAP ( A =>	FA3_l4_c49_Cout, B =>	FA2_l4_c49_Cout, CIN 	=>	FA1_l4_c49_Cout, S =>	FA1_l3_c50_S, COUT 	=>	FA1_l3_c50_Cout );

	FA2_l3_c50  : FA 
	PORT MAP ( A =>	FA3_l4_c50_S, B =>	FA2_l4_c50_S, CIN 	=>	FA1_l4_c50_S, S =>	FA2_l3_c50_S, COUT 	=>	FA2_l3_c50_Cout );

	FA1_l3_c51  : FA 
	PORT MAP ( A =>	FA3_l4_c50_Cout, B =>	FA2_l4_c50_Cout, CIN 	=>	FA1_l4_c50_Cout, S =>	FA1_l3_c51_S, COUT 	=>	FA1_l3_c51_Cout );

	FA2_l3_c51  : FA 
	PORT MAP ( A =>	FA3_l4_c51_S, B =>	FA2_l4_c51_S, CIN 	=>	FA1_l4_c51_S, S =>	FA2_l3_c51_S, COUT 	=>	FA2_l3_c51_Cout );

	FA1_l3_c52  : FA 
	PORT MAP ( A =>	FA3_l4_c51_Cout, B =>	FA2_l4_c51_Cout, CIN 	=>	FA1_l4_c51_Cout, S =>	FA1_l3_c52_S, COUT 	=>	FA1_l3_c52_Cout );

	FA2_l3_c52  : FA 
	PORT MAP ( A =>	HA1_l4_c52_S, B =>	FA2_l4_c52_S, CIN 	=>	FA1_l4_c52_S, S =>	FA2_l3_c52_S, COUT 	=>	FA2_l3_c52_Cout );

	FA1_l3_c53  : FA
	PORT MAP ( A =>	HA1_l4_c52_Cout, B =>	FA2_l4_c52_Cout, CIN 	=>	FA1_l4_c52_Cout, S =>	FA1_l3_c53_S, COUT 	=>	FA1_l3_c53_Cout );

	FA2_l3_c53  : FA 
	PORT MAP ( A =>	FA2_l4_c53_S, B =>	FA1_l4_c53_S, CIN 	=>	PP16(21), S =>	FA2_l3_c53_S, COUT 	=>	FA2_l3_c53_Cout );

	FA1_l3_c54  : FA 
	PORT MAP ( A =>	FA2_l4_c53_Cout, B =>	FA1_l4_c53_Cout, CIN 	=>	HA1_l4_c54_S, S =>	FA1_l3_c54_S, COUT 	=>	FA1_l3_c54_Cout );

	FA2_l3_c54  : FA 
	PORT MAP ( A =>	FA1_l4_c54_S, B =>	PP15(24), CIN 	=>	PP16(22), S =>	FA2_l3_c54_S, COUT 	=>	FA2_l3_c54_Cout );

	FA1_l3_c55  : FA 
	PORT MAP ( A =>	HA1_l4_c54_Cout, B =>	FA1_l4_c54_Cout, CIN 	=>	FA1_l4_c55_S, S =>	FA1_l3_c55_S, COUT 	=>	FA1_l3_c55_Cout );

	FA2_l3_c55  : FA 
	PORT MAP ( A =>	PP14(27), B =>	PP15(25), CIN 	=>	PP16(23), S =>	FA2_l3_c55_S, COUT 	=>	FA2_l3_c55_Cout );

	FA1_l3_c56  : FA 
	PORT MAP ( A =>	FA1_l4_c55_Cout, B =>	HA1_l4_c56_S, CIN 	=>	PP13(30), S =>	FA1_l3_c56_S, COUT 	=>	FA1_l3_c56_Cout );

	FA2_l3_c56  : FA 
	PORT MAP ( A =>	PP14(28), B =>	PP15(26), CIN 	=>	PP16(24), S =>	FA2_l3_c56_S, COUT 	=>	FA2_l3_c56_Cout );

	FA1_l3_c57  : FA 
	PORT MAP ( A =>	HA1_l4_c56_Cout, B =>	PP12_neg, CIN 	=>	PP13(31), S =>	FA1_l3_c57_S, COUT 	=>	FA1_l3_c57_Cout );

	FA2_l3_c57  : FA 
	PORT MAP ( A =>	PP14(29), B =>	PP15(27), CIN 	=>	PP16(25), S =>	FA2_l3_c57_S, COUT 	=>	FA2_l3_c57_Cout );

	FA1_l3_c58  : FA 
	PORT MAP ( A =>	'1', B =>	PP13(32), CIN 	=>	PP14(30), S =>	FA1_l3_c58_S, COUT 	=>	FA1_l3_c58_Cout );

	HA1_l3_c58  : HA 
	PORT MAP ( A =>	PP15(28), B =>	PP16(26), S =>	HA1_l3_c58_S, COUT 	=>	HA1_l3_c58_Cout );

	FA1_l3_c59  : FA 
	PORT MAP ( A =>	PP13_neg, B =>	PP14(31), CIN 	=>	PP15(29), S =>	FA1_l3_c59_S, COUT 	=>	FA1_l3_c59_Cout );

	HA1_l3_c60  : HA 
	PORT MAP ( A =>	'1', B =>	PP14(32), S =>	HA1_l3_c60_S, COUT 	=>	HA1_l3_c60_Cout );

	HA1_l2_c4  : HA 
	PORT MAP ( A =>	PP0(4), B =>	PP1(2), S =>	HA1_l2_c4_S, COUT 	=>	HA1_l2_c4_Cout );

	HA1_l2_c5  : HA 
	PORT MAP ( A =>	PP0(5), B =>	PP1(3), S =>	HA1_l2_c5_S, COUT 	=>	HA1_l2_c5_Cout );

	FA1_l2_c6  : FA 
	PORT MAP ( A =>	HA1_l3_c6_S, B =>	PP2(2), CIN 	=>	PP3(0), S =>	FA1_l2_c6_S, COUT 	=>	FA1_l2_c6_Cout );

	FA1_l2_c7  : FA 
	PORT MAP ( A =>	HA1_l3_c6_Cout, B =>	HA1_l3_c7_S, CIN 	=>	PP2(3), S =>	FA1_l2_c7_S, COUT 	=>	FA1_l2_c7_Cout );

	FA1_l2_c8  : FA 
	PORT MAP ( A =>	HA1_l3_c7_Cout, B =>	HA1_l3_c8_S, CIN 	=>	FA1_l3_c8_S, S =>	FA1_l2_c8_S, COUT 	=>	FA1_l2_c8_Cout );
	
	FA1_l2_c9  : FA 
	PORT MAP ( A =>	HA1_l3_c8_Cout, B =>	FA1_l3_c8_Cout, CIN 	=>	HA1_l3_c9_S, S =>	FA1_l2_c9_S, COUT 	=>	FA1_l2_c9_Cout );

	FA1_l2_c10  : FA 
	PORT MAP ( A =>	HA1_l3_c9_Cout, B =>	FA1_l3_c9_Cout, CIN 	=>	FA2_l3_c10_S, S =>	FA1_l2_c10_S, COUT 	=>	FA1_l2_c10_Cout );

	FA1_l2_c11  : FA 
	PORT MAP ( A =>	FA2_l3_c10_Cout, B =>	FA1_l3_c10_Cout, CIN 	=>	FA2_l3_c11_S, S =>	FA1_l2_c11_S, COUT 	=>	FA1_l2_c11_Cout );

	FA1_l2_c12  : FA 
	PORT MAP ( A =>	FA2_l3_c11_Cout, B =>	FA1_l3_c11_Cout, CIN 	=>	FA2_l3_c12_S, S =>	FA1_l2_c12_S, COUT 	=>	FA1_l2_c12_Cout );

	FA1_l2_c13  : FA 
	PORT MAP ( A =>	FA2_l3_c12_Cout, B =>	FA1_l3_c12_Cout, CIN 	=>	FA2_l3_c13_S, S =>	FA1_l2_c13_S, COUT 	=>	FA1_l2_c13_Cout );

	FA1_l2_c14  : FA 
	PORT MAP ( A =>	FA2_l3_c13_Cout, B =>	FA1_l3_c13_Cout, CIN 	=>	FA2_l3_c14_S, S =>	FA1_l2_c14_S, COUT 	=>	FA1_l2_c14_Cout );

	FA1_l2_c15  : FA
	PORT MAP ( A =>	FA2_l3_c14_Cout, B =>	FA1_l3_c14_Cout, CIN 	=>	FA2_l3_c15_S, S =>	FA1_l2_c15_S, COUT 	=>	FA1_l2_c15_Cout );

	FA1_l2_c16  : FA 
	PORT MAP ( A =>	FA2_l3_c15_Cout, B =>	FA1_l3_c15_Cout, CIN 	=>	FA2_l3_c16_S, S =>	FA1_l2_c16_S, COUT 	=>	FA1_l2_c16_Cout );

	FA1_l2_c17  : FA 
	PORT MAP ( A =>	FA2_l3_c16_Cout, B =>	FA1_l3_c16_Cout, CIN 	=>	FA2_l3_c17_S, S =>	FA1_l2_c17_S, COUT 	=>	FA1_l2_c17_Cout );

	FA1_l2_c18  : FA 
	PORT MAP ( A =>	FA2_l3_c17_Cout, B =>	FA1_l3_c17_Cout, CIN 	=>	FA2_l3_c18_S, S =>	FA1_l2_c18_S, COUT 	=>	FA1_l2_c18_Cout );

	FA1_l2_c19  : FA 
	PORT MAP ( A =>	FA2_l3_c18_Cout, B =>	FA1_l3_c18_Cout, CIN 	=>	FA2_l3_c19_S, S =>	FA1_l2_c19_S, COUT 	=>	FA1_l2_c19_Cout );

	FA1_l2_c20  : FA 
	PORT MAP ( A =>	FA2_l3_c19_Cout, B =>	FA1_l3_c19_Cout, CIN 	=>	FA2_l3_c20_S, S =>	FA1_l2_c20_S, COUT 	=>	FA1_l2_c20_Cout );

	FA1_l2_c21  : FA 
	PORT MAP ( A =>	FA2_l3_c20_Cout, B =>	FA1_l3_c20_Cout, CIN 	=>	FA2_l3_c21_S, S =>	FA1_l2_c21_S, COUT 	=>	FA1_l2_c21_Cout );

	FA1_l2_c22  : FA 
	PORT MAP ( A =>	FA2_l3_c21_Cout, B =>	FA1_l3_c21_Cout, CIN 	=>	FA2_l3_c22_S, S =>	FA1_l2_c22_S, COUT 	=>	FA1_l2_c22_Cout );

	FA1_l2_c23  : FA 
	PORT MAP ( A =>	FA2_l3_c22_Cout, B =>	FA1_l3_c22_Cout, CIN 	=>	FA2_l3_c23_S, S =>	FA1_l2_c23_S, COUT 	=>	FA1_l2_c23_Cout );

	FA1_l2_c24  : FA 
	PORT MAP ( A =>	FA2_l3_c23_Cout, B =>	FA1_l3_c23_Cout, CIN 	=>	FA2_l3_c24_S, S =>	FA1_l2_c24_S, COUT 	=>	FA1_l2_c24_Cout );

	FA1_l2_c25  : FA 
	PORT MAP ( A =>	FA2_l3_c24_Cout, B =>	FA1_l3_c24_Cout, CIN 	=>	FA2_l3_c25_S, S =>	FA1_l2_c25_S, COUT 	=>	FA1_l2_c25_Cout );

	FA1_l2_c26  : FA 
	PORT MAP ( A =>	FA2_l3_c25_Cout, B =>	FA1_l3_c25_Cout, CIN 	=>	FA2_l3_c26_S, S =>	FA1_l2_c26_S, COUT 	=>	FA1_l2_c26_Cout );

	FA1_l2_c27  : FA 
	PORT MAP ( A =>	FA2_l3_c26_Cout, B =>	FA1_l3_c26_Cout, CIN 	=>	FA2_l3_c27_S, S =>	FA1_l2_c27_S, COUT 	=>	FA1_l2_c27_Cout );

	FA1_l2_c28  : FA 
	PORT MAP ( A =>	FA2_l3_c27_Cout, B =>	FA1_l3_c27_Cout, CIN 	=>	FA2_l3_c28_S, S =>	FA1_l2_c28_S, COUT 	=>	FA1_l2_c28_Cout );

	FA1_l2_c29  : FA 
	PORT MAP ( A =>	FA2_l3_c28_Cout, B =>	FA1_l3_c28_Cout, CIN 	=>	FA2_l3_c29_S, S =>	FA1_l2_c29_S, COUT 	=>	FA1_l2_c29_Cout );

	FA1_l2_c30  : FA 
	PORT MAP ( A =>	FA2_l3_c29_Cout, B =>	FA1_l3_c29_Cout, CIN 	=>	FA2_l3_c30_S, S =>	FA1_l2_c30_S, COUT 	=>	FA1_l2_c30_Cout );

	FA1_l2_c31  : FA 
	PORT MAP ( A =>	FA2_l3_c30_Cout, B =>	FA1_l3_c30_Cout, CIN 	=>	FA2_l3_c31_S, S =>	FA1_l2_c31_S, COUT 	=>	FA1_l2_c31_Cout );

	FA1_l2_c32  : FA 
	PORT MAP ( A =>	FA2_l3_c31_Cout, B =>	FA1_l3_c31_Cout, CIN 	=>	FA2_l3_c32_S, S =>	FA1_l2_c32_S, COUT 	=>	FA1_l2_c32_Cout );

	FA1_l2_c33  : FA 
	PORT MAP ( A =>	FA2_l3_c32_Cout, B =>	FA1_l3_c32_Cout, CIN 	=>	FA2_l3_c33_S, S =>	FA1_l2_c33_S, COUT 	=>	FA1_l2_c33_Cout );

	FA1_l2_c34  : FA 
	PORT MAP ( A =>	FA2_l3_c33_Cout, B =>	FA1_l3_c33_Cout, CIN 	=>	FA2_l3_c34_S, S =>	FA1_l2_c34_S, COUT 	=>	FA1_l2_c34_Cout );

	FA1_l2_c35  : FA 
	PORT MAP ( A =>	FA2_l3_c34_Cout, B =>	FA1_l3_c34_Cout, CIN 	=>	FA2_l3_c35_S, S =>	FA1_l2_c35_S, COUT 	=>	FA1_l2_c35_Cout );

	FA1_l2_c36  : FA 
	PORT MAP ( A =>	FA2_l3_c35_Cout, B =>	FA1_l3_c35_Cout, CIN 	=>	FA2_l3_c36_S, S =>	FA1_l2_c36_S, COUT 	=>	FA1_l2_c36_Cout );

	FA1_l2_c37  : FA 
	PORT MAP ( A =>	FA2_l3_c36_Cout, B =>	FA1_l3_c36_Cout, CIN 	=>	FA2_l3_c37_S, S =>	FA1_l2_c37_S, COUT 	=>	FA1_l2_c37_Cout );

	FA1_l2_c38  : FA
	PORT MAP ( A =>	FA2_l3_c37_Cout, B =>	FA1_l3_c37_Cout, CIN 	=>	FA2_l3_c38_S, S =>	FA1_l2_c38_S, COUT 	=>	FA1_l2_c38_Cout );

	FA1_l2_c39  : FA 
	PORT MAP ( A =>	FA2_l3_c38_Cout, B =>	FA1_l3_c38_Cout, CIN 	=>	FA2_l3_c39_S, S =>	FA1_l2_c39_S, COUT 	=>	FA1_l2_c39_Cout );

	FA1_l2_c40  : FA 
	PORT MAP ( A =>	FA2_l3_c39_Cout, B =>	FA1_l3_c39_Cout, CIN 	=>	FA2_l3_c40_S, S =>	FA1_l2_c40_S, COUT 	=>	FA1_l2_c40_Cout );

	FA1_l2_c41  : FA 
	PORT MAP ( A =>	FA2_l3_c40_Cout, B =>	FA1_l3_c40_Cout, CIN 	=>	FA2_l3_c41_S, S =>	FA1_l2_c41_S, COUT 	=>	FA1_l2_c41_Cout );

	FA1_l2_c42  : FA 
	PORT MAP ( A =>	FA2_l3_c41_Cout, B =>	FA1_l3_c41_Cout, CIN 	=>	FA2_l3_c42_S, S =>	FA1_l2_c42_S, COUT 	=>	FA1_l2_c42_Cout );

	FA1_l2_c43  : FA 
	PORT MAP ( A =>	FA2_l3_c42_Cout, B =>	FA1_l3_c42_Cout, CIN 	=>	FA2_l3_c43_S, S =>	FA1_l2_c43_S, COUT 	=>	FA1_l2_c43_Cout );

	FA1_l2_c44  : FA 
	PORT MAP ( A =>	FA2_l3_c43_Cout, B =>	FA1_l3_c43_Cout, CIN 	=>	FA2_l3_c44_S, S =>	FA1_l2_c44_S, COUT 	=>	FA1_l2_c44_Cout );

	FA1_l2_c45  : FA 
	PORT MAP ( A =>	FA2_l3_c44_Cout, B =>	FA1_l3_c44_Cout, CIN 	=>	FA2_l3_c45_S, S =>	FA1_l2_c45_S, COUT 	=>	FA1_l2_c45_Cout );

	FA1_l2_c46  : FA 
	PORT MAP ( A =>	FA2_l3_c45_Cout, B =>	FA1_l3_c45_Cout, CIN 	=>	FA2_l3_c46_S, S =>	FA1_l2_c46_S, COUT 	=>	FA1_l2_c46_Cout );

	FA1_l2_c47  : FA 
	PORT MAP ( A =>	FA2_l3_c46_Cout, B =>	FA1_l3_c46_Cout, CIN 	=>	FA2_l3_c47_S, S =>	FA1_l2_c47_S, COUT 	=>	FA1_l2_c47_Cout );

	FA1_l2_c48  : FA 
	PORT MAP ( A =>	FA2_l3_c47_Cout, B =>	FA1_l3_c47_Cout, CIN 	=>	FA2_l3_c48_S, S =>	FA1_l2_c48_S, COUT 	=>	FA1_l2_c48_Cout );

	FA1_l2_c49  : FA 
	PORT MAP ( A =>	FA2_l3_c48_Cout, B =>	FA1_l3_c48_Cout, CIN 	=>	FA2_l3_c49_S, S =>	FA1_l2_c49_S, COUT 	=>	FA1_l2_c49_Cout );

	FA1_l2_c50  : FA 
	PORT MAP ( A =>	FA2_l3_c49_Cout, B =>	FA1_l3_c49_Cout, CIN 	=>	FA2_l3_c50_S, S =>	FA1_l2_c50_S, COUT 	=>	FA1_l2_c50_Cout );

	FA1_l2_c51  : FA 
	PORT MAP ( A =>	FA2_l3_c50_Cout, B =>	FA1_l3_c50_Cout, CIN 	=>	FA2_l3_c51_S, S =>	FA1_l2_c51_S, COUT 	=>	FA1_l2_c51_Cout );

	FA1_l2_c52  : FA 
	PORT MAP ( A =>	FA2_l3_c51_Cout, B =>	FA1_l3_c51_Cout, CIN 	=>	FA2_l3_c52_S, S =>	FA1_l2_c52_S, COUT 	=>	FA1_l2_c52_Cout );

	FA1_l2_c53  : FA 
	PORT MAP ( A =>	FA2_l3_c52_Cout, B =>	FA1_l3_c52_Cout, CIN 	=>	FA2_l3_c53_S, S =>	FA1_l2_c53_S, COUT 	=>	FA1_l2_c53_Cout );

	FA1_l2_c54  : FA 
	PORT MAP ( A =>	FA2_l3_c53_Cout, B =>	FA1_l3_c53_Cout, CIN 	=>	FA2_l3_c54_S, S =>	FA1_l2_c54_S, COUT 	=>	FA1_l2_c54_Cout );

	FA1_l2_c55  : FA 
	PORT MAP ( A =>	FA2_l3_c54_Cout, B =>	FA1_l3_c54_Cout, CIN 	=>	FA2_l3_c55_S, S =>	FA1_l2_c55_S, COUT 	=>	FA1_l2_c55_Cout );

	FA1_l2_c56  : FA 
	PORT MAP ( A =>	FA2_l3_c55_Cout, B =>	FA1_l3_c55_Cout, CIN 	=>	FA2_l3_c56_S, S =>	FA1_l2_c56_S, COUT 	=>	FA1_l2_c56_Cout );

	FA1_l2_c57  : FA 
	PORT MAP ( A =>	FA2_l3_c56_Cout, B =>	FA1_l3_c56_Cout, CIN 	=>	FA2_l3_c57_S, S =>	FA1_l2_c57_S, COUT 	=>	FA1_l2_c57_Cout );

	FA1_l2_c58  : FA 
	PORT MAP ( A =>	FA2_l3_c57_Cout, B =>	FA1_l3_c57_Cout, CIN 	=>	HA1_l3_c58_S, S =>	FA1_l2_c58_S, COUT 	=>	FA1_l2_c58_Cout );

	FA1_l2_c59  : FA 
	PORT MAP ( A =>	HA1_l3_c58_Cout, B =>	FA1_l3_c58_Cout, CIN 	=>	FA1_l3_c59_S, S =>	FA1_l2_c59_S, COUT 	=>	FA1_l2_c59_Cout );

	FA1_l2_c60  : FA 
	PORT MAP ( A =>	FA1_l3_c59_Cout, B =>	HA1_l3_c60_S, CIN 	=>	PP15(30), S =>	FA1_l2_c60_S, COUT 	=>	FA1_l2_c60_Cout );

	FA1_l2_c61  : FA 
	PORT MAP ( A =>	HA1_l3_c60_Cout, B =>	PP14_neg, CIN 	=>	PP15(31), S =>	FA1_l2_c61_S, COUT 	=>	FA1_l2_c61_Cout );

	HA1_l2_c62  : HA 
	PORT MAP ( A =>	'1', B =>	PP15(32), S =>	HA1_l2_c62_S, COUT 	=>	HA1_l2_c62_Cout );

	HA1_l1_c2  : HA 
	PORT MAP ( A =>	PP0(2), B =>	PP1(0), S =>	HA1_l1_c2_S, COUT 	=>	HA1_l1_c2_Cout );

	HA1_l1_c3  : HA 
	PORT MAP ( A =>	PP0(3), B =>	PP1(1), S =>	HA1_l1_c3_S, COUT 	=>	HA1_l1_c3_Cout );

	FA1_l1_c4  : FA 
	PORT MAP ( A =>	HA1_l2_c4_S, B =>	PP2(0), CIN 	=>	PP2(32), S =>	FA1_l1_c4_S, COUT 	=>	FA1_l1_c4_Cout );

	FA1_l1_c5  : FA 
	PORT MAP ( A =>	HA1_l2_c4_Cout, B =>	HA1_l2_c5_S, CIN 	=>	PP2(1), S =>	FA1_l1_c5_S, COUT 	=>	FA1_l1_c5_Cout );

	FA1_l1_c6  : FA 
	PORT MAP ( A =>	HA1_l2_c5_Cout, B =>	FA1_l2_c6_S, CIN 	=>	PP3(32), S =>	FA1_l1_c6_S, COUT 	=>	FA1_l1_c6_Cout );

	FA1_l1_c7  : FA
	PORT MAP ( A =>	FA1_l2_c6_Cout, B =>	FA1_l2_c7_S, CIN 	=>	PP3(1), S =>	FA1_l1_c7_S, COUT 	=>	FA1_l1_c7_Cout );

	FA1_l1_c8  : FA 
	PORT MAP ( A =>	FA1_l2_c7_Cout, B =>	FA1_l2_c8_S, CIN 	=>	PP4(32), S =>	FA1_l1_c8_S, COUT 	=>	FA1_l1_c8_Cout );

	FA1_l1_c9  : FA 
	PORT MAP ( A =>	FA1_l2_c8_Cout, B =>	FA1_l2_c9_S, CIN 	=>	FA1_l3_c9_S, S =>	FA1_l1_c9_S, COUT 	=>	FA1_l1_c9_Cout );

	FA1_l1_c10  : FA 
	PORT MAP ( A =>	FA1_l2_c9_Cout, B =>	FA1_l2_c10_S, CIN 	=>	FA1_l3_c10_S, S =>	FA1_l1_c10_S, COUT 	=>	FA1_l1_c10_Cout );

	FA1_l1_c11  : FA 
	PORT MAP ( A =>	FA1_l2_c10_Cout, B =>	FA1_l2_c11_S, CIN 	=>	FA1_l3_c11_S, S =>	FA1_l1_c11_S, COUT 	=>	FA1_l1_c11_Cout );

	FA1_l1_c12  : FA 
	PORT MAP ( A =>	FA1_l2_c11_Cout, B =>	FA1_l2_c12_S, CIN 	=>	FA1_l3_c12_S, S =>	FA1_l1_c12_S, COUT 	=>	FA1_l1_c12_Cout );

	FA1_l1_c13  : FA 
	PORT MAP ( A =>	FA1_l2_c12_Cout, B =>	FA1_l2_c13_S, CIN 	=>	FA1_l3_c13_S, S =>	FA1_l1_c13_S, COUT 	=>	FA1_l1_c13_Cout );

	FA1_l1_c14  : FA 
	PORT MAP ( A =>	FA1_l2_c13_Cout, B =>	FA1_l2_c14_S, CIN 	=>	FA1_l3_c14_S, S =>	FA1_l1_c14_S, COUT 	=>	FA1_l1_c14_Cout );

	FA1_l1_c15  : FA 
	PORT MAP ( A =>	FA1_l2_c14_Cout, B =>	FA1_l2_c15_S, CIN 	=>	FA1_l3_c15_S, S =>	FA1_l1_c15_S, COUT 	=>	FA1_l1_c15_Cout );

	FA1_l1_c16  : FA 
	PORT MAP ( A =>	FA1_l2_c15_Cout, B =>	FA1_l2_c16_S, CIN 	=>	FA1_l3_c16_S, S =>	FA1_l1_c16_S, COUT 	=>	FA1_l1_c16_Cout );

	FA1_l1_c17  : FA 
	PORT MAP ( A =>	FA1_l2_c16_Cout, B =>	FA1_l2_c17_S, CIN 	=>	FA1_l3_c17_S, S =>	FA1_l1_c17_S, COUT 	=>	FA1_l1_c17_Cout );

	FA1_l1_c18  : FA 
	PORT MAP ( A =>	FA1_l2_c17_Cout, B =>	FA1_l2_c18_S, CIN 	=>	FA1_l3_c18_S, S =>	FA1_l1_c18_S, COUT 	=>	FA1_l1_c18_Cout );

	FA1_l1_c19  : FA 
	PORT MAP ( A =>	FA1_l2_c18_Cout, B =>	FA1_l2_c19_S, CIN 	=>	FA1_l3_c19_S, S =>	FA1_l1_c19_S, COUT 	=>	FA1_l1_c19_Cout );

	FA1_l1_c20  : FA 
	PORT MAP ( A =>	FA1_l2_c19_Cout, B =>	FA1_l2_c20_S, CIN 	=>	FA1_l3_c20_S, S =>	FA1_l1_c20_S, COUT 	=>	FA1_l1_c20_Cout );

	FA1_l1_c21  : FA 
	PORT MAP ( A =>	FA1_l2_c20_Cout, B =>	FA1_l2_c21_S, CIN 	=>	FA1_l3_c21_S, S =>	FA1_l1_c21_S, COUT 	=>	FA1_l1_c21_Cout );

	FA1_l1_c22  : FA 
	PORT MAP ( A =>	FA1_l2_c21_Cout, B =>	FA1_l2_c22_S, CIN 	=>	FA1_l3_c22_S, S =>	FA1_l1_c22_S, COUT 	=>	FA1_l1_c22_Cout );

	FA1_l1_c23  : FA 
	PORT MAP ( A =>	FA1_l2_c22_Cout, B =>	FA1_l2_c23_S, CIN 	=>	FA1_l3_c23_S, S =>	FA1_l1_c23_S, COUT 	=>	FA1_l1_c23_Cout );

	FA1_l1_c24  : FA 
	PORT MAP ( A =>	FA1_l2_c23_Cout, B =>	FA1_l2_c24_S, CIN 	=>	FA1_l3_c24_S, S =>	FA1_l1_c24_S, COUT 	=>	FA1_l1_c24_Cout );

	FA1_l1_c25  : FA 
	PORT MAP ( A =>	FA1_l2_c24_Cout, B =>	FA1_l2_c25_S, CIN 	=>	FA1_l3_c25_S, S =>	FA1_l1_c25_S, COUT 	=>	FA1_l1_c25_Cout );

	FA1_l1_c26  : FA 
	PORT MAP ( A =>	FA1_l2_c25_Cout, B =>	FA1_l2_c26_S, CIN 	=>	FA1_l3_c26_S, S =>	FA1_l1_c26_S, COUT 	=>	FA1_l1_c26_Cout );

	FA1_l1_c27  : FA 
	PORT MAP ( A =>	FA1_l2_c26_Cout, B =>	FA1_l2_c27_S, CIN 	=>	FA1_l3_c27_S, S =>	FA1_l1_c27_S, COUT 	=>	FA1_l1_c27_Cout );

	FA1_l1_c28  : FA 
	PORT MAP ( A =>	FA1_l2_c27_Cout, B =>	FA1_l2_c28_S, CIN 	=>	FA1_l3_c28_S, S =>	FA1_l1_c28_S, COUT 	=>	FA1_l1_c28_Cout );

	FA1_l1_c29  : FA 
	PORT MAP ( A =>	FA1_l2_c28_Cout, B =>	FA1_l2_c29_S, CIN 	=>	FA1_l3_c29_S, S =>	FA1_l1_c29_S, COUT 	=>	FA1_l1_c29_Cout );

	FA1_l1_c30  : FA 
	PORT MAP ( A =>	FA1_l2_c29_Cout, B =>	FA1_l2_c30_S, CIN 	=>	FA1_l3_c30_S, S =>	FA1_l1_c30_S, COUT 	=>	FA1_l1_c30_Cout );

	FA1_l1_c31  : FA 
	PORT MAP ( A =>	FA1_l2_c30_Cout, B =>	FA1_l2_c31_S, CIN 	=>	FA1_l3_c31_S, S =>	FA1_l1_c31_S, COUT 	=>	FA1_l1_c31_Cout );

	FA1_l1_c32  : FA 
	PORT MAP ( A =>	FA1_l2_c31_Cout, B =>	FA1_l2_c32_S, CIN 	=>	FA1_l3_c32_S, S =>	FA1_l1_c32_S, COUT 	=>	FA1_l1_c32_Cout );

	FA1_l1_c33  : FA 
	PORT MAP ( A =>	FA1_l2_c32_Cout, B =>	FA1_l2_c33_S, CIN 	=>	FA1_l3_c33_S, S =>	FA1_l1_c33_S, COUT 	=>	FA1_l1_c33_Cout );

	FA1_l1_c34  : FA 
	PORT MAP ( A =>	FA1_l2_c33_Cout, B =>	FA1_l2_c34_S, CIN 	=>	FA1_l3_c34_S, S =>	FA1_l1_c34_S, COUT 	=>	FA1_l1_c34_Cout );

	FA1_l1_c35  : FA 
	PORT MAP ( A =>	FA1_l2_c34_Cout, B =>	FA1_l2_c35_S, CIN 	=>	FA1_l3_c35_S, S =>	FA1_l1_c35_S, COUT 	=>	FA1_l1_c35_Cout );

	FA1_l1_c36  : FA 
	PORT MAP ( A =>	FA1_l2_c35_Cout, B =>	FA1_l2_c36_S, CIN 	=>	FA1_l3_c36_S, S =>	FA1_l1_c36_S, COUT 	=>	FA1_l1_c36_Cout );

	FA1_l1_c37  : FA 
	PORT MAP ( A =>	FA1_l2_c36_Cout, B =>	FA1_l2_c37_S, CIN 	=>	FA1_l3_c37_S, S =>	FA1_l1_c37_S, COUT 	=>	FA1_l1_c37_Cout );

	FA1_l1_c38  : FA 
	PORT MAP ( A =>	FA1_l2_c37_Cout, B =>	FA1_l2_c38_S, CIN 	=>	FA1_l3_c38_S, S =>	FA1_l1_c38_S, COUT 	=>	FA1_l1_c38_Cout );

	FA1_l1_c39  : FA 
	PORT MAP ( A =>	FA1_l2_c38_Cout, B =>	FA1_l2_c39_S, CIN 	=>	FA1_l3_c39_S, S =>	FA1_l1_c39_S, COUT 	=>	FA1_l1_c39_Cout );

	FA1_l1_c40  : FA 
	PORT MAP ( A =>	FA1_l2_c39_Cout, B =>	FA1_l2_c40_S, CIN 	=>	FA1_l3_c40_S, S =>	FA1_l1_c40_S, COUT 	=>	FA1_l1_c40_Cout );

	FA1_l1_c41  : FA 
	PORT MAP ( A =>	FA1_l2_c40_Cout, B =>	FA1_l2_c41_S, CIN 	=>	FA1_l3_c41_S, S =>	FA1_l1_c41_S, COUT 	=>	FA1_l1_c41_Cout );

	FA1_l1_c42  : FA 
	PORT MAP ( A =>	FA1_l2_c41_Cout, B =>	FA1_l2_c42_S, CIN 	=>	FA1_l3_c42_S, S =>	FA1_l1_c42_S, COUT 	=>	FA1_l1_c42_Cout );

	FA1_l1_c43  : FA 
	PORT MAP ( A =>	FA1_l2_c42_Cout, B =>	FA1_l2_c43_S, CIN 	=>	FA1_l3_c43_S, S =>	FA1_l1_c43_S, COUT 	=>	FA1_l1_c43_Cout );

	FA1_l1_c44  : FA 
	PORT MAP ( A =>	FA1_l2_c43_Cout, B =>	FA1_l2_c44_S, CIN 	=>	FA1_l3_c44_S, S =>	FA1_l1_c44_S, COUT 	=>	FA1_l1_c44_Cout );

	FA1_l1_c45  : FA 
	PORT MAP ( A =>	FA1_l2_c44_Cout, B =>	FA1_l2_c45_S, CIN 	=>	FA1_l3_c45_S, S =>	FA1_l1_c45_S, COUT 	=>	FA1_l1_c45_Cout );

	FA1_l1_c46  : FA 
	PORT MAP ( A =>	FA1_l2_c45_Cout, B =>	FA1_l2_c46_S, CIN 	=>	FA1_l3_c46_S, S =>	FA1_l1_c46_S, COUT 	=>	FA1_l1_c46_Cout );

	FA1_l1_c47  : FA 
	PORT MAP ( A =>	FA1_l2_c46_Cout, B =>	FA1_l2_c47_S, CIN 	=>	FA1_l3_c47_S, S =>	FA1_l1_c47_S, COUT 	=>	FA1_l1_c47_Cout );

	FA1_l1_c48  : FA 
	PORT MAP ( A =>	FA1_l2_c47_Cout, B =>	FA1_l2_c48_S, CIN 	=>	FA1_l3_c48_S, S =>	FA1_l1_c48_S, COUT 	=>	FA1_l1_c48_Cout );

	FA1_l1_c49  : FA 
	PORT MAP ( A =>	FA1_l2_c48_Cout, B =>	FA1_l2_c49_S, CIN 	=>	FA1_l3_c49_S, S =>	FA1_l1_c49_S, COUT 	=>	FA1_l1_c49_Cout );

	FA1_l1_c50  : FA 
	PORT MAP ( A =>	FA1_l2_c49_Cout, B =>	FA1_l2_c50_S, CIN 	=>	FA1_l3_c50_S, S =>	FA1_l1_c50_S, COUT 	=>	FA1_l1_c50_Cout );

	FA1_l1_c51  : FA 
	PORT MAP ( A =>	FA1_l2_c50_Cout, B =>	FA1_l2_c51_S, CIN 	=>	FA1_l3_c51_S, S =>	FA1_l1_c51_S, COUT 	=>	FA1_l1_c51_Cout );

	FA1_l1_c52  : FA 
	PORT MAP ( A =>	FA1_l2_c51_Cout, B =>	FA1_l2_c52_S, CIN 	=>	FA1_l3_c52_S, S =>	FA1_l1_c52_S, COUT 	=>	FA1_l1_c52_Cout );

	FA1_l1_c53  : FA 
	PORT MAP ( A =>	FA1_l2_c52_Cout, B =>	FA1_l2_c53_S, CIN 	=>	FA1_l3_c53_S, S =>	FA1_l1_c53_S, COUT 	=>	FA1_l1_c53_Cout );

	FA1_l1_c54  : FA 
	PORT MAP ( A =>	FA1_l2_c53_Cout, B =>	FA1_l2_c54_S, CIN 	=>	FA1_l3_c54_S, S =>	FA1_l1_c54_S, COUT 	=>	FA1_l1_c54_Cout );

	FA1_l1_c55  : FA 
	PORT MAP ( A =>	FA1_l2_c54_Cout, B =>	FA1_l2_c55_S, CIN 	=>	FA1_l3_c55_S, S =>	FA1_l1_c55_S, COUT 	=>	FA1_l1_c55_Cout );

	FA1_l1_c56  : FA 
	PORT MAP ( A =>	FA1_l2_c55_Cout, B =>	FA1_l2_c56_S, CIN 	=>	FA1_l3_c56_S, S =>	FA1_l1_c56_S, COUT 	=>	FA1_l1_c56_Cout );

	FA1_l1_c57  : FA 
	PORT MAP ( A =>	FA1_l2_c56_Cout, B =>	FA1_l2_c57_S, CIN 	=>	FA1_l3_c57_S, S =>	FA1_l1_c57_S, COUT 	=>	FA1_l1_c57_Cout );

	FA1_l1_c58  : FA 
	PORT MAP ( A =>	FA1_l2_c57_Cout, B =>	FA1_l2_c58_S, CIN 	=>	FA1_l3_c58_S, S =>	FA1_l1_c58_S, COUT 	=>	FA1_l1_c58_Cout );

	FA1_l1_c59  : FA 
	PORT MAP ( A =>	FA1_l2_c58_Cout, B =>	FA1_l2_c59_S, CIN 	=>	PP16(27), S =>	FA1_l1_c59_S, COUT 	=>	FA1_l1_c59_Cout );

	FA1_l1_c60  : FA 
	PORT MAP ( A =>	FA1_l2_c59_Cout, B =>	FA1_l2_c60_S, CIN 	=>	PP16(28), S =>	FA1_l1_c60_S, COUT 	=>	FA1_l1_c60_Cout );

	FA1_l1_c61  : FA 
	PORT MAP ( A =>	FA1_l2_c60_Cout, B =>	FA1_l2_c61_S, CIN 	=>	PP16(29), S =>	FA1_l1_c61_S, COUT 	=>	FA1_l1_c61_Cout );

	FA1_l1_c62  : FA 
	PORT MAP ( A =>	FA1_l2_c61_Cout, B =>	HA1_l2_c62_S, CIN 	=>	PP16(30), S =>	FA1_l1_c62_S, COUT 	=>	FA1_l1_c62_Cout );

	FA1_l1_c63  : FA 
	PORT MAP ( A =>	HA1_l2_c62_Cout, B =>	PP15_neg, CIN 	=>	PP16(31), S =>	FA1_l1_c63_S, COUT 	=>	FA1_l1_c63_Cout ); 
	
	---- last sum ----
	process (sum_1,sum_2)
	
	begin  
		
		sum <= unsigned(sum_1) + unsigned(sum_2);
		M <= std_logic_vector(sum);
	
	end process;

end behavior;
